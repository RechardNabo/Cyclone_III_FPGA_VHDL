-- ============================================================================
-- 2-to-1 Multiplexer Implementation - Programming Guidance
-- ============================================================================
-- 
-- PROJECT OVERVIEW:
-- This file implements a 2-to-1 Multiplexer (MUX), which is a fundamental
-- digital circuit that selects one of two input signals based on a select
-- control signal. The multiplexer routes the selected input to the output,
-- making it essential for data routing, signal switching, and conditional
-- data flow in digital systems.
--
-- LEARNING OBJECTIVES:
-- 1. Understand multiplexer operation and selection logic
-- 2. Learn conditional signal routing in VHDL
-- 3. Practice control signal implementation
-- 4. Explore data path design fundamentals
--
-- ============================================================================
-- STEP-BY-STEP IMPLEMENTATION GUIDE:
-- ============================================================================
--
-- STEP 1: LIBRARY DECLARATIONS
-- ----------------------------------------------------------------------------
-- Required Libraries:
-- - IEEE library for standard logic types
-- - std_logic_1164 package for std_logic and logical operators
-- - numeric_std package for arithmetic operations (optional)
-- 
-- TODO: Add library IEEE;
-- TODO: Add use IEEE.std_logic_1164.all;
-- TODO: Add use IEEE.numeric_std.all; (for advanced implementations)
--
-- ============================================================================
-- STEP 2: ENTITY DECLARATION
-- ----------------------------------------------------------------------------
-- The entity defines the 2-to-1 multiplexer interface
--
-- Entity Requirements:
-- - Name: mux_2to1 (maintain current naming convention)
-- - Inputs: I0, I1 (two data inputs), S (select signal)
-- - Output: Y (selected output)
-- - All signals are single-bit std_logic
--
-- Port Specifications:
-- - I0 : in std_logic (Data input 0)
-- - I1 : in std_logic (Data input 1)
-- - S  : in std_logic (Select signal)
-- - Y  : out std_logic (Output)
--
-- TODO: Declare entity with appropriate port map
-- TODO: Add port comments for clarity
-- TODO: Consider signal naming conventions
--
-- ============================================================================
-- STEP 3: ARCHITECTURE IMPLEMENTATION
-- ============================================================================
-- Multiple approaches to implement 2-to-1 multiplexer functionality:
--
-- OPTION A: BEHAVIORAL MODELING (Process-based)
-- - Use process with complete sensitivity list
-- - Implement with if-else or case statements
-- - Good for understanding selection logic
-- - Easy to extend and modify
--
-- OPTION B: DATAFLOW MODELING (Concurrent assignments)
-- - Use Boolean expressions for output
-- - Direct implementation of selection logic
-- - Most efficient and clear approach
-- - Excellent synthesis results
--
-- OPTION C: CONDITIONAL ASSIGNMENTS
-- - Use when-else statements for output
-- - Clear conditional logic representation
-- - Good for understanding input-output relationships
--
-- OPTION D: SELECTED ASSIGNMENTS
-- - Use with-select statements
-- - Compact truth table representation
-- - Good for systematic implementation
--
-- OPTION E: STRUCTURAL MODELING
-- - Use basic gates (AND, OR, NOT)
-- - Demonstrates gate-level implementation
-- - Good for understanding hardware structure
-- - Educational value for logic design
--
-- ============================================================================
-- 2-TO-1 MULTIPLEXER TRUTH TABLE:
-- ============================================================================
--
-- Inputs     | Output
-- I1  I0  S  | Y     | Description
-- -----------|-------|----------------------------------
-- 0   0   0  | 0     | Select I0 (0)
-- 0   1   0  | 1     | Select I0 (1)
-- 1   0   0  | 0     | Select I0 (0)
-- 1   1   0  | 1     | Select I0 (1)
-- 0   0   1  | 0     | Select I1 (0)
-- 0   1   1  | 0     | Select I1 (0)
-- 1   0   1  | 1     | Select I1 (1)
-- 1   1   1  | 1     | Select I1 (1)
--
-- Simplified Truth Table:
-- S | Y
-- --|--------
-- 0 | I0
-- 1 | I1
--
-- Key Insights:
-- - When S = 0, output Y = I0
-- - When S = 1, output Y = I1
-- - Select signal controls which input passes through
-- - Non-selected input is ignored
--
-- ============================================================================
-- IMPLEMENTATION CONSIDERATIONS:
-- ============================================================================
--
-- BOOLEAN EXPRESSIONS:
-- Output Expression:
-- - Y = S'·I0 + S·I1 (Sum of products form)
-- - Y = S ? I1 : I0 (Conditional expression)
-- - Y = (NOT S AND I0) OR (S AND I1)
--
-- GATE-LEVEL IMPLEMENTATION:
-- - Two AND gates for input selection
-- - One OR gate for output combination
-- - One NOT gate for select inversion
-- - Total: 4 gates for complete implementation
--
-- VHDL IMPLEMENTATION TECHNIQUES:
-- - Use 'when-else' for conditional assignment
-- - Use 'with-select' for systematic selection
-- - Use Boolean expression for direct implementation
-- - Use process with if-else for behavioral modeling
--
-- SYNTHESIS CONSIDERATIONS:
-- - Multiplexer maps efficiently to FPGA LUT resources
-- - Typically requires 1 LUT for 2-to-1 MUX
-- - Very efficient resource utilization
-- - Synthesis tools optimize automatically
--
-- TIMING CHARACTERISTICS:
-- - Propagation delay from inputs to output
-- - Select signal has critical timing path
-- - Consider setup and hold times for all inputs
-- - Glitch-free operation important for data integrity
--
-- ============================================================================
-- 2-TO-1 MULTIPLEXER APPLICATIONS:
-- ============================================================================
--
-- 1. DATA ROUTING AND SWITCHING:
--    - Route data between different sources
--    - Switch between alternate data paths
--    - Implement data selectors in processors
--    - Create configurable data connections
--
-- 2. CONDITIONAL DATA FLOW:
--    - Select between different computational results
--    - Implement conditional assignments
--    - Create decision-making circuits
--    - Control data flow based on conditions
--
-- 3. BUILDING LARGER MULTIPLEXERS:
--    - Combine multiple 2-to-1 MUX to create 4-to-1, 8-to-1, etc.
--    - Hierarchical multiplexer design
--    - Tree structure for large multiplexers
--    - Scalable multiplexer architectures
--
-- 4. PROCESSOR DESIGN:
--    - ALU input selection
--    - Register file output selection
--    - Instruction decode logic
--    - Control unit implementation
--
-- 5. MEMORY SYSTEMS:
--    - Address multiplexing
--    - Data path selection
--    - Memory bank selection
--    - Cache line selection
--
-- 6. COMMUNICATION SYSTEMS:
--    - Channel selection
--    - Protocol switching
--    - Data stream multiplexing
--    - Signal routing matrices
--
-- 7. CONTROL LOGIC:
--    - Mode selection circuits
--    - Configuration switching
--    - State-dependent routing
--    - Conditional control paths
--
-- ============================================================================
-- TESTING STRATEGY:
-- ============================================================================
--
-- BASIC FUNCTIONALITY TESTS:
-- 1. Test Case 1: S=0, I0=0, I1=X → Expected: Y=0
-- 2. Test Case 2: S=0, I0=1, I1=X → Expected: Y=1
-- 3. Test Case 3: S=1, I0=X, I1=0 → Expected: Y=0
-- 4. Test Case 4: S=1, I0=X, I1=1 → Expected: Y=1
--
-- SELECTION VERIFICATION:
-- - Verify correct input selection for S=0 (I0 selected)
-- - Verify correct input selection for S=1 (I1 selected)
-- - Test with all combinations of I0 and I1 values
-- - Confirm non-selected input doesn't affect output
--
-- BOOLEAN LOGIC VERIFICATION:
-- - Confirm Boolean expression: Y = S'·I0 + S·I1
-- - Test with all 8 possible input combinations
-- - Verify truth table compliance
-- - Check for unexpected output states
--
-- TIMING ANALYSIS:
-- - Measure propagation delays from all inputs
-- - Verify setup and hold time requirements
-- - Test for glitches during select transitions
-- - Validate simultaneous input changes
--
-- METAVALUE HANDLING:
-- - Test with 'X' (unknown) inputs → Expected behavior
-- - Test with 'Z' (high-impedance) inputs → Expected behavior
-- - Test with 'U' (uninitialized) inputs → Expected behavior
-- - Verify proper metavalue propagation
--
-- EDGE CASE TESTING:
-- - Rapid select signal transitions
-- - Simultaneous input and select changes
-- - Hold time violations
-- - Setup time violations
--
-- ============================================================================
-- RECOMMENDED IMPLEMENTATION APPROACH:
-- ============================================================================
--
-- FOR BEGINNERS:
-- 1. Start with truth table analysis and understanding
-- 2. Implement using when-else conditional assignment
-- 3. Create comprehensive testbench covering all cases
-- 4. Understand selection logic operation
--
-- FOR INTERMEDIATE USERS:
-- 1. Implement multiple architectures (behavioral, dataflow)
-- 2. Compare synthesis results between approaches
-- 3. Analyze timing characteristics
-- 4. Create structural implementation using basic gates
--
-- FOR ADVANCED USERS:
-- 1. Use 2-to-1 MUX as component in larger multiplexers
-- 2. Create parameterized multi-bit multiplexer
-- 3. Optimize for specific FPGA architectures
-- 4. Implement advanced routing structures
--
-- ============================================================================
-- EXTENSION EXERCISES:
-- ============================================================================
--
-- 1. MULTI-BIT 2-TO-1 MULTIPLEXER:
--    - Create N-bit 2-to-1 multiplexer for vector inputs
--    - Use generate statements for scalability
--    - Implement bus-width parameterization
--    - Compare with individual bit multiplexers
--
-- 2. 4-TO-1 MULTIPLEXER FROM 2-TO-1:
--    - Create 4-to-1 MUX using three 2-to-1 MUX
--    - Understand hierarchical design methodology
--    - Compare with direct 4-to-1 implementation
--    - Analyze resource utilization differences
--
-- 3. 8-TO-1 MULTIPLEXER TREE:
--    - Build 8-to-1 MUX using 2-to-1 building blocks
--    - Implement tree structure design
--    - Create scalable multiplexer architecture
--    - Add parameterization for different sizes
--
-- 4. TRI-STATE MULTIPLEXER:
--    - Add enable signal for tri-state output
--    - Implement high-impedance state control
--    - Create bus-compatible multiplexer
--    - Add output enable functionality
--
-- 5. MULTIPLEXER WITH PRIORITY:
--    - Implement priority-based selection
--    - Add multiple select signals
--    - Create priority encoder integration
--    - Implement conflict resolution logic
--
-- 6. GLITCH-FREE MULTIPLEXER:
--    - Implement break-before-make switching
--    - Add delay elements for glitch prevention
--    - Create clean switching transitions
--    - Analyze timing requirements
--
-- ============================================================================
-- COMMON MISTAKES TO AVOID:
-- ============================================================================
--
-- 1. INCORRECT SELECTION LOGIC:
--    - Don't confuse select signal polarity
--    - Ensure correct input-to-output mapping
--    - Verify selection logic against truth table
--    - Test all selection combinations thoroughly
--
-- 2. SENSITIVITY LIST ERRORS:
--    - Include all input signals in process sensitivity list
--    - Missing signals cause simulation/synthesis mismatch
--    - Use 'all' keyword for automatic sensitivity (VHDL-2008)
--    - Avoid incomplete sensitivity lists
--
-- 3. SIGNAL ASSIGNMENT ISSUES:
--    - Use concurrent assignments for combinational logic
--    - Avoid creating unintended latches
--    - Ensure output is always assigned
--    - Don't mix clocked and combinational logic
--
-- 4. TIMING CONSIDERATIONS:
--    - Consider propagation delays through selection logic
--    - Account for select signal timing requirements
--    - Avoid glitches during select transitions
--    - Understand critical path timing
--
-- 5. METAVALUE HANDLING:
--    - Properly handle unknown select signals
--    - Define behavior for undefined inputs
--    - Consider initialization requirements
--    - Test with realistic signal conditions
--
-- ============================================================================
-- DESIGN VERIFICATION CHECKLIST:
-- ============================================================================
--
-- □ Entity declaration includes all input and output ports
-- □ Port directions correctly specified (in/out)
-- □ All 8 input combinations tested exhaustively
-- □ Selection logic verified (S=0 selects I0, S=1 selects I1)
-- □ Boolean expression matches truth table
-- □ No undefined or uninitialized output states
-- □ Metavalue behavior tested and understood
-- □ Synthesis completes without errors or warnings
-- □ Timing requirements satisfied
-- □ Resource utilization acceptable
-- □ Code follows project VHDL style guidelines
-- □ Comments clearly explain multiplexer functionality
-- □ Testbench provides complete coverage
-- □ Glitch-free operation verified
--
-- ============================================================================
-- MULTIPLEXER IN DIGITAL DESIGN CONTEXT:
-- ============================================================================
--
-- RELATIONSHIP TO OTHER CIRCUITS:
-- - Building block for larger multiplexers
-- - Component in data path design
-- - Used in control logic implementation
-- - Foundation for routing networks
--
-- BOOLEAN ALGEBRA PROPERTIES:
-- - Demonstrates conditional logic principles
-- - Illustrates sum-of-products implementation
-- - Shows gate-level design methodology
-- - Foundation for understanding selection logic
--
-- DATA PATH DESIGN:
-- - Essential component in processor design
-- - Used for register file implementation
-- - Critical in ALU input selection
-- - Important for memory addressing
--
-- ============================================================================
-- PHYSICAL IMPLEMENTATION NOTES:
-- ============================================================================
--
-- FPGA IMPLEMENTATION:
-- - Typically uses 1 LUT for 2-to-1 multiplexer
-- - Very efficient resource utilization
-- - Can be implemented in single logic element
-- - Modern FPGAs optimize automatically
--
-- TIMING CHARACTERISTICS:
-- - tpd_sel: Propagation delay from select to output
-- - tpd_data: Propagation delay from data inputs to output
-- - tsu: Setup time for input signals
-- - th: Hold time for input signals
-- - Consider select signal critical path
--
-- POWER CONSUMPTION:
-- - Static: Minimal leakage current
-- - Dynamic: Switching power depends on activity
-- - Select signal transitions affect power most
-- - Input switching power varies with selection
--
-- GLITCH CONSIDERATIONS:
-- - Select signal changes can cause output glitches
-- - Input transitions during selection can cause glitches
-- - Consider glitch-free design for critical applications
-- - Use synchronous design to minimize glitches
--
-- ============================================================================
-- ADVANCED MULTIPLEXER CONCEPTS:
-- ============================================================================
--
-- HIERARCHICAL DESIGN:
-- - Use 2-to-1 MUX to build larger multiplexers
-- - Tree structure for N-to-1 multiplexers
-- - Logarithmic delay scaling with size
-- - Modular design approach
--
-- TRANSMISSION GATE IMPLEMENTATION:
-- - CMOS transmission gate multiplexers
-- - Bidirectional signal flow capability
-- - Lower propagation delay
-- - Reduced power consumption
--
-- MULTIPLEXER NETWORKS:
-- - Crossbar switch implementation
-- - Routing fabric in FPGAs
-- - Network-on-chip routing
-- - Interconnection networks
--
-- OPTIMIZATION TECHNIQUES:
-- - Select signal buffering for large fan-out
-- - Pipeline registers for high-speed operation
-- - Parallel multiplexer structures
-- - Custom layout for performance
--
-- ============================================================================
-- SIMULATION AND VERIFICATION NOTES:
-- ============================================================================
--
-- TESTBENCH REQUIREMENTS:
-- - Exhaustive testing of all 8 input combinations
-- - Selection logic verification
-- - Boolean expression verification
-- - Timing analysis with appropriate delays
--
-- WAVEFORM ANALYSIS:
-- - Verify correct input selection behavior
-- - Check for glitches during select transitions
-- - Validate propagation delay characteristics
-- - Confirm proper initialization behavior
--
-- COVERAGE ANALYSIS:
-- - Functional coverage for all input combinations
-- - Toggle coverage for all input and output signals
-- - Path coverage for both selection paths
-- - Assertion coverage for selection properties
--
-- FORMAL VERIFICATION:
-- - Prove selection correctness: Y = S ? I1 : I0
-- - Verify Boolean expression equivalence
-- - Check truth table compliance
-- - Validate timing constraints and requirements
--
-- ASSERTION-BASED VERIFICATION:
-- - Assert correct selection behavior
-- - Check for proper output assignment
-- - Verify no undefined output states
-- - Validate timing relationships
--
-- ============================================================================
-- COMPARISON WITH OTHER MULTIPLEXERS:
-- ============================================================================
--
-- 2-TO-1 vs 4-TO-1 MULTIPLEXER:
-- - 2-to-1: 1 select bit, simpler logic
-- - 4-to-1: 2 select bits, more complex
-- - 2-to-1 more efficient for binary selection
-- - 4-to-1 better for multiple option selection
--
-- RESOURCE COMPARISON:
-- - 2-to-1 MUX: 1 LUT, minimal resources
-- - 4-to-1 MUX: 1 LUT, same resources in FPGA
-- - Larger MUX: Multiple LUTs, tree structure
-- - Choice depends on application requirements
--
-- PERFORMANCE COMPARISON:
-- - 2-to-1 MUX: Minimal propagation delay
-- - Larger MUX: Logarithmic delay increase
-- - Tree structure affects timing
-- - Consider critical path requirements
--
-- ============================================================================
-- MULTIPLEXER DESIGN PATTERNS:
-- ============================================================================
--
-- BASIC SELECTION PATTERN:
-- - Simple input selection based on control
-- - Most common multiplexer usage
-- - Direct implementation of selection logic
-- - Suitable for most applications
--
-- HIERARCHICAL PATTERN:
-- - Build larger MUX from smaller ones
-- - Modular and scalable design
-- - Easy to understand and maintain
-- - Good for complex routing requirements
--
-- PARAMETERIZED PATTERN:
-- - Generic multiplexer with configurable size
-- - Use generics for width and select bits
-- - Reusable component design
-- - Suitable for library development
--
-- PIPELINE PATTERN:
-- - Add registers for high-speed operation
-- - Break critical paths with flip-flops
-- - Increase throughput at cost of latency
-- - Suitable for high-frequency designs
--
-- ============================================================================
-- IMPLEMENTATION TEMPLATE:
-- ============================================================================
--
-- [Add your library declarations here]
--
-- [Add your entity declaration here]
--
-- [Add your architecture implementation here]
--
-- ============================================================================