-- ============================================================================
-- N-Bit Parameterized Counter Implementation - Programming Guidance
-- ============================================================================
-- 
-- PROJECT OVERVIEW:
-- This file implements a parameterized N-bit binary counter that can be
-- configured for any bit width. This generic design provides flexibility
-- for different applications while maintaining consistent functionality.
-- The counter supports various counting modes, control signals, and can
-- be easily scaled from small 4-bit counters to large 32-bit or wider
-- counters for different system requirements.
--
-- LEARNING OBJECTIVES:
-- 1. Understand VHDL generic parameters and parameterized design
-- 2. Learn scalable sequential logic implementation
-- 3. Practice generic type conversions and calculations
-- 4. Explore resource optimization for different bit widths
-- 5. Understand parameterized testbench development
--
-- ============================================================================
-- STEP-BY-STEP IMPLEMENTATION GUIDE:
-- ============================================================================
--
-- STEP 1: LIBRARY DECLARATIONS
-- ----------------------------------------------------------------------------
-- Required Libraries:
-- - IEEE library for standard logic types
-- - std_logic_1164 package for std_logic and logical operators
-- - numeric_std package for arithmetic operations (strongly recommended)
-- - math_real package for mathematical functions (for generic calculations)
-- 
-- TODO: Add library IEEE;
-- TODO: Add use IEEE.std_logic_1164.all;
-- TODO: Add use IEEE.numeric_std.all;
-- TODO: Add use IEEE.math_real.all; (for log2 calculations)
--
-- ============================================================================
-- STEP 2: ENTITY DECLARATION WITH GENERICS
-- ============================================================================
-- The entity defines the parameterized interface for the N-bit counter
--
-- Generic Parameters:
-- - N : positive := 8 (Default bit width, must be positive)
-- - RESET_VALUE : natural := 0 (Default reset value)
-- - COUNT_UP : boolean := true (Default count direction)
-- - ASYNC_RESET : boolean := true (Reset type selection)
--
-- Entity Requirements:
-- - Name: counter_nbit (maintain current naming convention)
-- - Generic parameters for configurability
-- - Inputs: Clock, reset, enable, load, direction control
-- - Outputs: N-bit count value, terminal count flags
-- - Scalable port definitions using generics
--
-- Port Specifications:
-- - clk : in std_logic (Clock input for synchronous operation)
-- - reset : in std_logic (Reset signal - async or sync based on generic)
-- - enable : in std_logic (Count enable control)
-- - load : in std_logic (Parallel load control)
-- - up_down : in std_logic (Count direction: '1' = up, '0' = down)
-- - load_data : in std_logic_vector(N-1 downto 0) (Parallel load data)
-- - count : out std_logic_vector(N-1 downto 0) (Current count value)
-- - tc_up : out std_logic (Terminal count up flag)
-- - tc_down : out std_logic (Terminal count down flag)
-- - carry_out : out std_logic (Carry output for cascading)
-- - borrow_out : out std_logic (Borrow output for cascading)
-- - overflow : out std_logic (Overflow detection flag)
-- - underflow : out std_logic (Underflow detection flag)
--
-- Generic Considerations:
-- - Bit width validation (N > 0)
-- - Reset value range checking (0 <= RESET_VALUE < 2^N)
-- - Default parameter selection
-- - Synthesis optimization hints
--
-- TODO: Declare entity with generic parameters
-- TODO: Add comprehensive port comments
-- TODO: Validate generic parameter ranges
-- TODO: Plan for maximum bit width support
--
-- ============================================================================
-- STEP 3: PARAMETERIZED COUNTER OPERATION DEFINITIONS
-- ============================================================================
--
-- PARAMETERIZED COUNTER PRINCIPLES:
-- - Scalable bit width from 1 to 32+ bits
-- - Generic-based terminal count calculation
-- - Configurable reset value and behavior
-- - Automatic overflow/underflow detection
-- - Resource optimization based on bit width
--
-- COUNTING RANGES:
-- - N-bit counter: 0 to (2^N - 1)
-- - 4-bit: 0 to 15
-- - 8-bit: 0 to 255
-- - 16-bit: 0 to 65535
-- - 32-bit: 0 to 4294967295
--
-- TERMINAL COUNT CALCULATIONS:
-- - MAX_COUNT = (2^N) - 1
-- - MIN_COUNT = 0
-- - TC_UP when count = MAX_COUNT
-- - TC_DOWN when count = MIN_COUNT
-- - Overflow when count wraps from MAX to 0
-- - Underflow when count wraps from 0 to MAX
--
-- GENERIC PARAMETER USAGE:
-- - Bit width: std_logic_vector(N-1 downto 0)
-- - Maximum value: (2**N) - 1
-- - Reset value: to_unsigned(RESET_VALUE, N)
-- - Type conversions: unsigned ↔ std_logic_vector
--
-- RESOURCE SCALING:
-- - Logic elements scale linearly with N
-- - Arithmetic resources increase with bit width
-- - Routing complexity grows with N
-- - Clock frequency may decrease with larger N
--
-- TODO: Calculate terminal count values using generics
-- TODO: Implement parameterized type conversions
-- TODO: Plan resource optimization strategies
-- TODO: Design overflow/underflow detection
--
-- ============================================================================
-- STEP 4: PARAMETERIZED ARCHITECTURE IMPLEMENTATION
-- ============================================================================
--
-- OPTION 1: GENERIC SYNCHRONOUS ARCHITECTURE
-- ----------------------------------------------------------------------------
-- Scalable synchronous counter with configurable parameters
--
-- Implementation Approach:
-- - Use generics for all size-dependent calculations
-- - Implement configurable reset behavior
-- - Support both synchronous and asynchronous reset
-- - Optimize for different bit widths
--
-- Example Structure:
-- architecture behavioral of counter_nbit is
--     -- Constants derived from generics
--     constant MAX_COUNT : unsigned(N-1 downto 0) := (others => '1');
--     constant MIN_COUNT : unsigned(N-1 downto 0) := (others => '0');
--     constant RESET_VAL : unsigned(N-1 downto 0) := to_unsigned(RESET_VALUE, N);
--     
--     -- Internal signals
--     signal count_reg : unsigned(N-1 downto 0) := RESET_VAL;
--     signal next_count : unsigned(N-1 downto 0);
--     
-- begin
--     -- Next count calculation
--     next_count_proc: process(count_reg, enable, up_down, load, load_data)
--     begin
--         if load = '1' then
--             next_count <= unsigned(load_data);
--         elsif enable = '1' then
--             if up_down = '1' then
--                 if count_reg = MAX_COUNT then
--                     next_count <= MIN_COUNT; -- Wraparound
--                 else
--                     next_count <= count_reg + 1;
--                 end if;
--             else
--                 if count_reg = MIN_COUNT then
--                     next_count <= MAX_COUNT; -- Wraparound
--                 else
--                     next_count <= count_reg - 1;
--                 end if;
--             end if;
--         else
--             next_count <= count_reg; -- Hold
--         end if;
--     end process;
--     
--     -- Clocked process (configurable reset type)
--     clocked_proc: process(clk, reset)
--     begin
--         if ASYNC_RESET and reset = '1' then
--             count_reg <= RESET_VAL;
--         elsif rising_edge(clk) then
--             if not ASYNC_RESET and reset = '1' then
--                 count_reg <= RESET_VAL;
--             else
--                 count_reg <= next_count;
--             end if;
--         end if;
--     end process;
--     
--     -- Output assignments
--     count <= std_logic_vector(count_reg);
--     tc_up <= '1' when count_reg = MAX_COUNT else '0';
--     tc_down <= '1' when count_reg = MIN_COUNT else '0';
--     overflow <= '1' when (count_reg = MAX_COUNT and enable = '1' and up_down = '1') else '0';
--     underflow <= '1' when (count_reg = MIN_COUNT and enable = '1' and up_down = '0') else '0';
--     carry_out <= tc_up and enable and up_down;
--     borrow_out <= tc_down and enable and not up_down;
-- end behavioral;
--
-- TODO: Implement generic constant calculations
-- TODO: Add configurable reset type support
-- TODO: Implement parameterized arithmetic operations
-- TODO: Generate appropriate terminal count flags
--
-- OPTION 2: OPTIMIZED SMALL COUNTER ARCHITECTURE
-- ----------------------------------------------------------------------------
-- Optimized implementation for small bit widths (N <= 8)
--
-- Implementation Approach:
-- - Use integer type for small counters
-- - Simplified arithmetic operations
-- - Reduced type conversion overhead
-- - Optimized for speed and area
--
-- Example Structure:
-- architecture optimized_small of counter_nbit is
--     signal count_int : integer range 0 to (2**N)-1 := RESET_VALUE;
--     constant MAX_VAL : integer := (2**N) - 1;
-- begin
--     counter_proc: process(clk, reset)
--     begin
--         if ASYNC_RESET and reset = '1' then
--             count_int <= RESET_VALUE;
--         elsif rising_edge(clk) then
--             if not ASYNC_RESET and reset = '1' then
--                 count_int <= RESET_VALUE;
--             elsif load = '1' then
--                 count_int <= to_integer(unsigned(load_data));
--             elsif enable = '1' then
--                 if up_down = '1' then
--                     if count_int = MAX_VAL then
--                         count_int <= 0;
--                     else
--                         count_int <= count_int + 1;
--                     end if;
--                 else
--                     if count_int = 0 then
--                         count_int <= MAX_VAL;
--                     else
--                         count_int <= count_int - 1;
--                     end if;
--                 end if;
--             end if;
--         end if;
--     end process;
--     
--     count <= std_logic_vector(to_unsigned(count_int, N));
--     tc_up <= '1' when count_int = MAX_VAL else '0';
--     tc_down <= '1' when count_int = 0 else '0';
-- end optimized_small;
--
-- TODO: Implement integer-based counting for small N
-- TODO: Add range constraints for integer signals
-- TODO: Optimize type conversions
-- TODO: Verify synthesis results for different N values
--
-- OPTION 3: LARGE COUNTER ARCHITECTURE
-- ----------------------------------------------------------------------------
-- Optimized implementation for large bit widths (N > 16)
--
-- Implementation Approach:
-- - Pipeline arithmetic operations for high frequency
-- - Separate increment/decrement logic
-- - Optimized carry chain implementation
-- - Resource balancing for large bit widths
--
-- Example Structure:
-- architecture large_counter of counter_nbit is
--     signal count_reg : unsigned(N-1 downto 0) := to_unsigned(RESET_VALUE, N);
--     signal increment : std_logic;
--     signal decrement : std_logic;
--     
--     -- Pipeline registers for large counters
--     signal count_pipe : unsigned(N-1 downto 0);
--     
-- begin
--     -- Control signal generation
--     increment <= enable and up_down and not load;
--     decrement <= enable and not up_down and not load;
--     
--     -- Pipelined counter for large bit widths
--     large_counter_proc: process(clk, reset)
--     begin
--         if ASYNC_RESET and reset = '1' then
--             count_reg <= to_unsigned(RESET_VALUE, N);
--             count_pipe <= to_unsigned(RESET_VALUE, N);
--         elsif rising_edge(clk) then
--             if not ASYNC_RESET and reset = '1' then
--                 count_reg <= to_unsigned(RESET_VALUE, N);
--                 count_pipe <= to_unsigned(RESET_VALUE, N);
--             else
--                 -- Pipeline stage 1: Prepare next value
--                 if load = '1' then
--                     count_pipe <= unsigned(load_data);
--                 elsif increment = '1' then
--                     count_pipe <= count_reg + 1;
--                 elsif decrement = '1' then
--                     count_pipe <= count_reg - 1;
--                 else
--                     count_pipe <= count_reg;
--                 end if;
--                 
--                 -- Pipeline stage 2: Update register
--                 count_reg <= count_pipe;
--             end if;
--         end if;
--     end process;
-- end large_counter;
--
-- TODO: Implement pipelined architecture for large N
-- TODO: Add carry chain optimization
-- TODO: Balance pipeline stages for timing
-- TODO: Verify timing closure for large bit widths
--
-- ============================================================================
-- STEP 5: ADVANCED PARAMETERIZED FEATURES
-- ============================================================================
--
-- CONFIGURABLE MODULUS COUNTER:
-- - Generic modulus parameter
-- - Runtime modulus configuration
-- - Automatic terminal count adjustment
-- - Flexible counting ranges
--
-- MULTI-MODE PARAMETERIZED COUNTER:
-- - Selectable counting modes via generics
-- - Binary, BCD, Gray code support
-- - Mode-specific optimizations
-- - Unified parameterized interface
--
-- CASCADABLE PARAMETERIZED COUNTER:
-- - Generic cascade width configuration
-- - Automatic carry/borrow chain generation
-- - Hierarchical counter structures
-- - Scalable multi-level counting
--
-- PERFORMANCE-OPTIMIZED COUNTER:
-- - Bit-width specific optimizations
-- - Synthesis directive integration
-- - FPGA-specific resource utilization
-- - Timing-driven implementation selection
--
-- FAULT-TOLERANT PARAMETERIZED COUNTER:
-- - Error detection and correction
-- - Redundant counting logic
-- - Parameterized reliability features
-- - Graceful degradation modes
--
-- TODO: Select appropriate advanced features
-- TODO: Implement parameterized enhancements
-- TODO: Add generic-based optimizations
-- TODO: Verify scalability across bit widths
--
-- ============================================================================
-- IMPLEMENTATION CONSIDERATIONS:
-- ============================================================================
--
-- GENERIC PARAMETER VALIDATION:
-- - Bit width range checking (1 <= N <= 32)
-- - Reset value validation (0 <= RESET_VALUE < 2^N)
-- - Boolean parameter consistency
-- - Synthesis tool compatibility
-- - Default parameter selection
--
-- PARAMETERIZED TYPE HANDLING:
-- - Generic-based vector sizing
-- - Dynamic type conversions
-- - Range constraint calculations
-- - Overflow/underflow detection
-- - Cross-bit-width compatibility
--
-- SYNTHESIS OPTIMIZATION:
-- - Bit-width specific optimizations
-- - Resource utilization balancing
-- - Timing constraint scaling
-- - Power optimization strategies
-- - FPGA architecture targeting
--
-- TESTABILITY CONSIDERATIONS:
-- - Parameterized testbench development
-- - Generic-based test pattern generation
-- - Scalable verification methodology
-- - Cross-bit-width testing
-- - Performance characterization
--
-- DOCUMENTATION REQUIREMENTS:
-- - Generic parameter descriptions
-- - Bit-width scaling guidelines
-- - Performance characteristics
-- - Resource utilization data
-- - Application examples
--
-- ============================================================================
-- APPLICATIONS:
-- ============================================================================
--
-- 1. SCALABLE TIMING SYSTEMS:
--    - Configurable timer bit widths
--    - Application-specific timing ranges
--    - Resource-optimized implementations
--    - Multi-resolution timing
--
-- 2. PARAMETERIZED ADDRESS GENERATION:
--    - Memory size-specific addressing
--    - Configurable address ranges
--    - Multi-level memory hierarchies
--    - Scalable DMA controllers
--
-- 3. FLEXIBLE FREQUENCY DIVISION:
--    - Configurable division ratios
--    - Multi-rate clock generation
--    - Scalable prescaler chains
--    - Application-specific frequencies
--
-- 4. CONFIGURABLE PROTOCOL COUNTERS:
--    - Protocol-specific bit widths
--    - Scalable packet counters
--    - Flexible sequence numbering
--    - Multi-protocol support
--
-- 5. PARAMETERIZED SIGNAL PROCESSING:
--    - Configurable sample counters
--    - Scalable buffer addressing
--    - Multi-rate processing
--    - Flexible window sizing
--
-- ============================================================================
-- TESTING STRATEGY:
-- ============================================================================
--
-- PARAMETERIZED FUNCTIONAL TESTING:
-- - Test multiple bit widths (4, 8, 16, 32)
-- - Verify generic parameter effects
-- - Cross-bit-width consistency
-- - Boundary condition testing
-- - Terminal count verification
--
-- GENERIC PARAMETER TESTING:
-- - Valid parameter range testing
-- - Invalid parameter handling
-- - Default parameter verification
-- - Parameter interaction testing
-- - Synthesis compatibility testing
--
-- SCALABILITY TESTING:
-- - Performance vs bit width analysis
-- - Resource utilization scaling
-- - Timing closure verification
-- - Power consumption characterization
-- - Maximum bit width determination
--
-- CROSS-CONFIGURATION TESTING:
-- - Different reset types
-- - Various counting modes
-- - Multiple modulus values
-- - Different default values
-- - Boolean parameter combinations
--
-- INTEGRATION TESTING:
-- - Multi-instance integration
-- - Cascaded counter chains
-- - System-level performance
-- - Cross-bit-width interfacing
-- - Real-world application testing
--
-- ============================================================================
-- RECOMMENDED IMPLEMENTATION APPROACH:
-- ============================================================================
--
-- FOR BEGINNERS:
-- 1. Start with simple 8-bit parameterized counter
-- 2. Add basic generic parameters (N, RESET_VALUE)
-- 3. Implement synchronous reset version
-- 4. Create parameterized testbench
-- 5. Test with different bit widths (4, 8, 16)
--
-- FOR INTERMEDIATE USERS:
-- 1. Add configurable reset type (sync/async)
-- 2. Implement advanced control features
-- 3. Add overflow/underflow detection
-- 4. Create comprehensive parameterized testbench
-- 5. Analyze resource scaling characteristics
--
-- FOR ADVANCED USERS:
-- 1. Implement bit-width specific optimizations
-- 2. Add performance-oriented architectures
-- 3. Create hierarchical parameterized design
-- 4. Implement advanced verification methodology
-- 5. Optimize for specific FPGA architectures
--
-- ============================================================================
-- EXTENSION EXERCISES:
-- ============================================================================
--
-- 1. MULTI-DIMENSIONAL PARAMETERIZED COUNTER:
--    - Multiple generic parameters
--    - Complex parameter relationships
--    - Multi-mode operation selection
--    - Advanced configuration options
--
-- 2. SELF-CONFIGURING COUNTER:
--    - Runtime parameter adjustment
--    - Dynamic bit width modification
--    - Adaptive performance optimization
--    - Intelligent resource allocation
--
-- 3. HIERARCHICAL PARAMETERIZED DESIGN:
--    - Multi-level counter structures
--    - Parameterized component instantiation
--    - Scalable system architectures
--    - Complex parameter propagation
--
-- 4. PERFORMANCE-ADAPTIVE COUNTER:
--    - Automatic architecture selection
--    - Bit-width specific optimizations
--    - Dynamic performance tuning
--    - Resource-aware implementation
--
-- 5. VERIFICATION-CENTRIC DESIGN:
--    - Built-in parameterized verification
--    - Self-testing capabilities
--    - Automated parameter validation
--    - Comprehensive coverage analysis
--
-- ============================================================================
-- COMMON MISTAKES TO AVOID:
-- ============================================================================
--
-- 1. GENERIC PARAMETER ISSUES:
--    - Invalid parameter ranges
--    - Inconsistent parameter usage
--    - Missing parameter validation
--    - Poor default parameter selection
--
-- 2. TYPE CONVERSION ERRORS:
--    - Incorrect generic-based sizing
--    - Type mismatch in assignments
--    - Range constraint violations
--    - Synthesis tool incompatibilities
--
-- 3. SCALABILITY PROBLEMS:
--    - Non-scalable implementation approaches
--    - Bit-width specific hardcoding
--    - Resource utilization inefficiencies
--    - Timing closure failures for large N
--
-- 4. TESTBENCH LIMITATIONS:
--    - Non-parameterized test patterns
--    - Insufficient bit-width coverage
--    - Missing generic parameter testing
--    - Inadequate scalability verification
--
-- 5. DOCUMENTATION DEFICIENCIES:
--    - Missing generic parameter descriptions
--    - Incomplete scaling guidelines
--    - Insufficient application examples
--    - Poor parameter interaction documentation
--
-- ============================================================================
-- DESIGN VERIFICATION CHECKLIST:
-- ============================================================================
--
-- □ Generic parameters properly declared and validated
-- □ Entity ports correctly sized using generics
-- □ All bit-width dependent calculations use generics
-- □ Type conversions handle all bit widths correctly
-- □ Terminal count calculations scale properly
-- □ Reset behavior consistent across bit widths
-- □ Synthesis results scale appropriately
-- □ Testbench parameterized for multiple bit widths
-- □ Documentation covers all generic parameters
-- □ Performance characterized across bit widths
-- □ Resource utilization analyzed and optimized
-- □ Timing closure verified for target bit widths
-- □ Cross-bit-width compatibility verified
-- □ Default parameters provide reasonable behavior
-- □ Error handling covers invalid parameters
--
-- ============================================================================
-- PHYSICAL IMPLEMENTATION NOTES:
-- ============================================================================
--
-- FPGA RESOURCE SCALING:
-- - Logic Elements: ~N LUTs for N-bit counter
-- - Registers: N flip-flops for count storage
-- - Routing: Increases with bit width
-- - Carry Chains: Utilized for arithmetic operations
-- - Clock Resources: Global clock distribution
--
-- BIT-WIDTH PERFORMANCE CHARACTERISTICS:
-- - 4-bit: ~500MHz, minimal resources
-- - 8-bit: ~400MHz, moderate resources
-- - 16-bit: ~300MHz, significant resources
-- - 32-bit: ~200MHz, substantial resources
-- - 64-bit: ~150MHz, extensive resources
--
-- OPTIMIZATION STRATEGIES:
-- - Small counters (N<=8): Use integer types
-- - Medium counters (8<N<=16): Standard unsigned
-- - Large counters (N>16): Consider pipelining
-- - Very large (N>32): Hierarchical approach
--
-- ============================================================================
-- IMPLEMENTATION TEMPLATE:
-- ============================================================================
--
-- [Add your library declarations here]
--
-- [Add your entity declaration with generics here]
--
-- [Add your parameterized architecture implementation here]
--
-- ============================================================================