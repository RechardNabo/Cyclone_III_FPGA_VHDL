-- ============================================================================
-- 4-to-1 Multiplexer Implementation - Programming Guidance
-- ============================================================================
-- 
-- PROJECT OVERVIEW:
-- This file implements a 4-to-1 Multiplexer (MUX), which is a digital circuit
-- that selects one of four input signals based on a 2-bit select control signal.
-- The multiplexer routes the selected input to the output, making it essential
-- for data routing, signal switching, and conditional data flow in larger
-- digital systems. This is an extension of the 2-to-1 multiplexer concept.
--
-- LEARNING OBJECTIVES:
-- 1. Understand multi-input multiplexer operation and selection logic
-- 2. Learn multi-bit control signal implementation in VHDL
-- 3. Practice hierarchical design using smaller multiplexers
-- 4. Explore scalable data path design fundamentals
--
-- ============================================================================
-- STEP-BY-STEP IMPLEMENTATION GUIDE:
-- ============================================================================
--
-- STEP 1: LIBRARY DECLARATIONS
-- ----------------------------------------------------------------------------
-- Required Libraries:
-- - IEEE library for standard logic types
-- - std_logic_1164 package for std_logic and logical operators
-- - numeric_std package for arithmetic operations (optional)
-- 
-- TODO: Add library IEEE;
-- TODO: Add use IEEE.std_logic_1164.all;
-- TODO: Add use IEEE.numeric_std.all; (for advanced implementations)
--
-- ============================================================================
-- STEP 2: ENTITY DECLARATION
-- ----------------------------------------------------------------------------
-- The entity defines the 4-to-1 multiplexer interface
--
-- Entity Requirements:
-- - Name: mux_4to1 (maintain current naming convention)
-- - Inputs: I0, I1, I2, I3 (four data inputs), S (2-bit select signal)
-- - Output: Y (selected output)
-- - Data signals are single-bit std_logic
-- - Select signal is 2-bit std_logic_vector
--
-- Port Specifications:
-- - I0 : in std_logic (Data input 0)
-- - I1 : in std_logic (Data input 1)
-- - I2 : in std_logic (Data input 2)
-- - I3 : in std_logic (Data input 3)
-- - S  : in std_logic_vector(1 downto 0) (2-bit select signal)
-- - Y  : out std_logic (Output)
--
-- TODO: Declare entity with appropriate port map
-- TODO: Add port comments for clarity
-- TODO: Consider signal naming conventions
--
-- ============================================================================
-- STEP 3: ARCHITECTURE IMPLEMENTATION
-- ============================================================================
-- Multiple approaches to implement 4-to-1 multiplexer functionality:
--
-- OPTION A: BEHAVIORAL MODELING (Process-based)
-- - Use process with complete sensitivity list
-- - Implement with case statement for select signal
-- - Good for understanding selection logic
-- - Easy to extend and modify
--
-- OPTION B: DATAFLOW MODELING (Concurrent assignments)
-- - Use Boolean expressions for output
-- - Direct implementation of selection logic
-- - Most efficient and clear approach
-- - Excellent synthesis results
--
-- OPTION C: CONDITIONAL ASSIGNMENTS
-- - Use when-else statements for output
-- - Clear conditional logic representation
-- - Good for understanding input-output relationships
--
-- OPTION D: SELECTED ASSIGNMENTS
-- - Use with-select statements
-- - Compact truth table representation
-- - Good for systematic implementation
--
-- OPTION E: STRUCTURAL MODELING
-- - Use three 2-to-1 multiplexers
-- - Demonstrates hierarchical design
-- - Good for understanding modular construction
-- - Educational value for scalable design
--
-- OPTION F: GATE-LEVEL IMPLEMENTATION
-- - Use basic gates (AND, OR, NOT)
-- - Demonstrates complete gate-level design
-- - Good for understanding hardware structure
-- - Educational value for logic design
--
-- ============================================================================
-- 4-TO-1 MULTIPLEXER TRUTH TABLE:
-- ============================================================================
--
-- Inputs        | Output
-- I3 I2 I1 I0 S | Y     | Description
-- --------------|-------|----------------------------------
-- X  X  X  0  00| 0     | Select I0 (0)
-- X  X  X  1  00| 1     | Select I0 (1)
-- X  X  0  X  01| 0     | Select I1 (0)
-- X  X  1  X  01| 1     | Select I1 (1)
-- X  0  X  X  10| 0     | Select I2 (0)
-- X  1  X  X  10| 1     | Select I2 (1)
-- 0  X  X  X  11| 0     | Select I3 (0)
-- 1  X  X  X  11| 1     | Select I3 (1)
--
-- Simplified Truth Table:
-- S[1:0] | Y
-- -------|--------
-- 00     | I0
-- 01     | I1
-- 10     | I2
-- 11     | I3
--
-- Key Insights:
-- - S = "00" selects I0
-- - S = "01" selects I1
-- - S = "10" selects I2
-- - S = "11" selects I3
-- - 2-bit select signal allows 4 input selection
-- - Non-selected inputs are ignored
--
-- ============================================================================
-- IMPLEMENTATION CONSIDERATIONS:
-- ============================================================================
--
-- BOOLEAN EXPRESSIONS:
-- Output Expression (Sum of Products):
-- - Y = S1'·S0'·I0 + S1'·S0·I1 + S1·S0'·I2 + S1·S0·I3
-- - Where S1 = S(1) and S0 = S(0)
--
-- HIERARCHICAL IMPLEMENTATION:
-- - First level: Two 2-to-1 MUX (I0,I1 and I2,I3)
-- - Second level: One 2-to-1 MUX (combines first level outputs)
-- - S(0) controls first level selection
-- - S(1) controls second level selection
--
-- GATE-LEVEL IMPLEMENTATION:
-- - Four AND gates for input selection (4 inputs each)
-- - One OR gate for output combination (4 inputs)
-- - Two NOT gates for select signal inversion
-- - Total: 7 gates for complete implementation
--
-- VHDL IMPLEMENTATION TECHNIQUES:
-- - Use 'case' statement for systematic selection
-- - Use 'when-else' for conditional assignment
-- - Use Boolean expression for direct implementation
-- - Use component instantiation for structural design
--
-- SYNTHESIS CONSIDERATIONS:
-- - 4-to-1 multiplexer maps efficiently to FPGA LUT resources
-- - Typically requires 1 LUT for 4-to-1 MUX
-- - Very efficient resource utilization
-- - Synthesis tools optimize automatically
--
-- TIMING CHARACTERISTICS:
-- - Propagation delay from inputs to output
-- - Select signal has critical timing path
-- - Consider setup and hold times for all inputs
-- - Decode delay for 2-bit select signal
--
-- ============================================================================
-- 4-TO-1 MULTIPLEXER APPLICATIONS:
-- ============================================================================
--
-- 1. DATA ROUTING AND SWITCHING:
--    - Route data between multiple sources
--    - Switch between four alternate data paths
--    - Implement data selectors in processors
--    - Create configurable data connections
--
-- 2. PROCESSOR DESIGN:
--    - ALU operand selection (4 sources)
--    - Register file output selection
--    - Instruction decode logic
--    - Control unit implementation
--    - Pipeline stage input selection
--
-- 3. MEMORY SYSTEMS:
--    - Memory bank selection (4 banks)
--    - Cache line selection
--    - Address multiplexing
--    - Data path selection
--    - Memory controller interfaces
--
-- 4. COMMUNICATION SYSTEMS:
--    - Channel selection (4 channels)
--    - Protocol switching
--    - Data stream multiplexing
--    - Signal routing matrices
--    - Interface selection
--
-- 5. CONTROL LOGIC:
--    - Mode selection circuits (4 modes)
--    - Configuration switching
--    - State-dependent routing
--    - Conditional control paths
--    - Function selection
--
-- 6. BUILDING LARGER MULTIPLEXERS:
--    - Combine multiple 4-to-1 MUX to create 8-to-1, 16-to-1, etc.
--    - Hierarchical multiplexer design
--    - Tree structure for large multiplexers
--    - Scalable multiplexer architectures
--
-- 7. DIGITAL SIGNAL PROCESSING:
--    - Input source selection for DSP algorithms
--    - Filter coefficient selection
--    - Data path configuration
--    - Algorithm mode selection
--
-- ============================================================================
-- TESTING STRATEGY:
-- ============================================================================
--
-- BASIC FUNCTIONALITY TESTS:
-- 1. Test Case 1: S="00", I0=0, I1=X, I2=X, I3=X → Expected: Y=0
-- 2. Test Case 2: S="00", I0=1, I1=X, I2=X, I3=X → Expected: Y=1
-- 3. Test Case 3: S="01", I0=X, I1=0, I2=X, I3=X → Expected: Y=0
-- 4. Test Case 4: S="01", I0=X, I1=1, I2=X, I3=X → Expected: Y=1
-- 5. Test Case 5: S="10", I0=X, I1=X, I2=0, I3=X → Expected: Y=0
-- 6. Test Case 6: S="10", I0=X, I1=X, I2=1, I3=X → Expected: Y=1
-- 7. Test Case 7: S="11", I0=X, I1=X, I2=X, I3=0 → Expected: Y=0
-- 8. Test Case 8: S="11", I0=X, I1=X, I2=X, I3=1 → Expected: Y=1
--
-- SELECTION VERIFICATION:
-- - Verify correct input selection for each S value
-- - Test with all combinations of input values
-- - Confirm non-selected inputs don't affect output
-- - Validate 2-bit select signal decoding
--
-- BOOLEAN LOGIC VERIFICATION:
-- - Confirm Boolean expression implementation
-- - Test with all 64 possible input combinations (4 data + 2 select)
-- - Verify truth table compliance
-- - Check for unexpected output states
--
-- TIMING ANALYSIS:
-- - Measure propagation delays from all inputs
-- - Verify setup and hold time requirements
-- - Test for glitches during select transitions
-- - Validate simultaneous input changes
-- - Check select signal decode timing
--
-- METAVALUE HANDLING:
-- - Test with 'X' (unknown) inputs → Expected behavior
-- - Test with 'Z' (high-impedance) inputs → Expected behavior
-- - Test with 'U' (uninitialized) inputs → Expected behavior
-- - Verify proper metavalue propagation
--
-- EDGE CASE TESTING:
-- - Rapid select signal transitions
-- - Simultaneous input and select changes
-- - Invalid select signal combinations (if applicable)
-- - Hold time violations
-- - Setup time violations
--
-- ============================================================================
-- RECOMMENDED IMPLEMENTATION APPROACH:
-- ============================================================================
--
-- FOR BEGINNERS:
-- 1. Start with truth table analysis and understanding
-- 2. Implement using case statement in process
-- 3. Create comprehensive testbench covering all cases
-- 4. Understand 2-bit select signal decoding
--
-- FOR INTERMEDIATE USERS:
-- 1. Implement multiple architectures (behavioral, dataflow)
-- 2. Compare synthesis results between approaches
-- 3. Analyze timing characteristics
-- 4. Create structural implementation using 2-to-1 MUX
--
-- FOR ADVANCED USERS:
-- 1. Use 4-to-1 MUX as component in larger multiplexers
-- 2. Create parameterized multi-bit multiplexer
-- 3. Optimize for specific FPGA architectures
-- 4. Implement advanced routing structures
--
-- ============================================================================
-- EXTENSION EXERCISES:
-- ============================================================================
--
-- 1. MULTI-BIT 4-TO-1 MULTIPLEXER:
--    - Create N-bit 4-to-1 multiplexer for vector inputs
--    - Use generate statements for scalability
--    - Implement bus-width parameterization
--    - Compare with individual bit multiplexers
--
-- 2. 8-TO-1 MULTIPLEXER FROM 4-TO-1:
--    - Create 8-to-1 MUX using two 4-to-1 MUX and one 2-to-1 MUX
--    - Understand hierarchical design methodology
--    - Compare with direct 8-to-1 implementation
--    - Analyze resource utilization differences
--
-- 3. 16-TO-1 MULTIPLEXER TREE:
--    - Build 16-to-1 MUX using 4-to-1 building blocks
--    - Implement tree structure design
--    - Create scalable multiplexer architecture
--    - Add parameterization for different sizes
--
-- 4. TRI-STATE 4-TO-1 MULTIPLEXER:
--    - Add enable signal for tri-state output
--    - Implement high-impedance state control
--    - Create bus-compatible multiplexer
--    - Add output enable functionality
--
-- 5. PRIORITY 4-TO-1 MULTIPLEXER:
--    - Implement priority-based selection
--    - Add priority encoder integration
--    - Create conflict resolution logic
--    - Handle multiple active inputs
--
-- 6. REGISTERED 4-TO-1 MULTIPLEXER:
--    - Add input and output registers
--    - Implement pipelined operation
--    - Create synchronous multiplexer
--    - Add clock and reset signals
--
-- ============================================================================
-- COMMON MISTAKES TO AVOID:
-- ============================================================================
--
-- 1. INCORRECT SELECTION LOGIC:
--    - Don't confuse select signal bit ordering
--    - Ensure correct input-to-output mapping
--    - Verify selection logic against truth table
--    - Test all selection combinations thoroughly
--
-- 2. SELECT SIGNAL HANDLING:
--    - Properly handle 2-bit select signal
--    - Use correct indexing for select bits
--    - Avoid confusion between S(1) and S(0)
--    - Consider select signal as std_logic_vector
--
-- 3. SENSITIVITY LIST ERRORS:
--    - Include all input signals in process sensitivity list
--    - Include complete select signal vector
--    - Missing signals cause simulation/synthesis mismatch
--    - Use 'all' keyword for automatic sensitivity (VHDL-2008)
--
-- 4. SIGNAL ASSIGNMENT ISSUES:
--    - Use concurrent assignments for combinational logic
--    - Avoid creating unintended latches
--    - Ensure output is always assigned
--    - Don't mix clocked and combinational logic
--
-- 5. CASE STATEMENT COMPLETENESS:
--    - Cover all possible select signal values
--    - Use 'others' clause for safety
--    - Avoid incomplete case statements
--    - Handle unexpected select values
--
-- 6. TIMING CONSIDERATIONS:
--    - Consider propagation delays through selection logic
--    - Account for select signal decode timing
--    - Avoid glitches during select transitions
--    - Understand critical path timing
--
-- ============================================================================
-- DESIGN VERIFICATION CHECKLIST:
-- ============================================================================
--
-- □ Entity declaration includes all input and output ports
-- □ Port directions correctly specified (in/out)
-- □ Select signal properly declared as std_logic_vector
-- □ All 16 selection combinations tested (4 select × 4 cases each)
-- □ Selection logic verified for each select value
-- □ Boolean expression matches truth table
-- □ No undefined or uninitialized output states
-- □ Case statement covers all select possibilities
-- □ 'Others' clause included for safety
-- □ Metavalue behavior tested and understood
-- □ Synthesis completes without errors or warnings
-- □ Timing requirements satisfied
-- □ Resource utilization acceptable
-- □ Code follows project VHDL style guidelines
-- □ Comments clearly explain multiplexer functionality
-- □ Testbench provides complete coverage
-- □ Glitch-free operation verified
--
-- ============================================================================
-- MULTIPLEXER IN DIGITAL DESIGN CONTEXT:
-- ============================================================================
--
-- RELATIONSHIP TO OTHER CIRCUITS:
-- - Building block for larger multiplexers
-- - Component in data path design
-- - Used in control logic implementation
-- - Foundation for routing networks
-- - Essential in processor design
--
-- BOOLEAN ALGEBRA PROPERTIES:
-- - Demonstrates multi-input selection logic
-- - Illustrates sum-of-products implementation
-- - Shows gate-level design methodology
-- - Foundation for understanding complex selection
--
-- DATA PATH DESIGN:
-- - Critical component in processor design
-- - Used for register file implementation
-- - Essential in ALU input selection
-- - Important for memory addressing
-- - Key in pipeline stage design
--
-- HIERARCHICAL DESIGN PRINCIPLES:
-- - Can be built from smaller multiplexers
-- - Demonstrates modular design approach
-- - Shows scalability concepts
-- - Illustrates design reuse principles
--
-- ============================================================================
-- PHYSICAL IMPLEMENTATION NOTES:
-- ============================================================================
--
-- FPGA IMPLEMENTATION:
-- - Typically uses 1 LUT for 4-to-1 multiplexer
-- - Very efficient resource utilization
-- - Can be implemented in single logic element
-- - Modern FPGAs optimize automatically
-- - LUT6 can handle 4-to-1 MUX easily
--
-- TIMING CHARACTERISTICS:
-- - tpd_sel: Propagation delay from select to output
-- - tpd_data: Propagation delay from data inputs to output
-- - tsu: Setup time for input signals
-- - th: Hold time for input signals
-- - tdecode: Select signal decode time
-- - Consider select signal critical path
--
-- POWER CONSUMPTION:
-- - Static: Minimal leakage current
-- - Dynamic: Switching power depends on activity
-- - Select signal transitions affect power most
-- - Input switching power varies with selection
-- - More inputs mean potentially higher power
--
-- GLITCH CONSIDERATIONS:
-- - Select signal changes can cause output glitches
-- - Input transitions during selection can cause glitches
-- - 2-bit select decode can create timing skew
-- - Consider glitch-free design for critical applications
-- - Use synchronous design to minimize glitches
--
-- ============================================================================
-- ADVANCED MULTIPLEXER CONCEPTS:
-- ============================================================================
--
-- HIERARCHICAL DESIGN:
-- - Use 2-to-1 MUX to build 4-to-1 MUX
-- - Tree structure for larger multiplexers
-- - Logarithmic delay scaling with size
-- - Modular design approach
-- - Design reuse benefits
--
-- TRANSMISSION GATE IMPLEMENTATION:
-- - CMOS transmission gate multiplexers
-- - Bidirectional signal flow capability
-- - Lower propagation delay
-- - Reduced power consumption
-- - Better analog signal handling
--
-- MULTIPLEXER NETWORKS:
-- - Crossbar switch implementation
-- - Routing fabric in FPGAs
-- - Network-on-chip routing
-- - Interconnection networks
-- - Matrix switching systems
--
-- OPTIMIZATION TECHNIQUES:
-- - Select signal buffering for large fan-out
-- - Pipeline registers for high-speed operation
-- - Parallel multiplexer structures
-- - Custom layout for performance
-- - Power optimization strategies
--
-- ============================================================================
-- SIMULATION AND VERIFICATION NOTES:
-- ============================================================================
--
-- TESTBENCH REQUIREMENTS:
-- - Exhaustive testing of all input combinations
-- - Selection logic verification for each select value
-- - Boolean expression verification
-- - Timing analysis with appropriate delays
-- - Edge case testing
--
-- WAVEFORM ANALYSIS:
-- - Verify correct input selection behavior
-- - Check for glitches during select transitions
-- - Validate propagation delay characteristics
-- - Confirm proper initialization behavior
-- - Analyze select signal decode timing
--
-- COVERAGE ANALYSIS:
-- - Functional coverage for all input combinations
-- - Toggle coverage for all input and output signals
-- - Path coverage for all selection paths
-- - Assertion coverage for selection properties
-- - State coverage for select signal values
--
-- FORMAL VERIFICATION:
-- - Prove selection correctness for each select value
-- - Verify Boolean expression equivalence
-- - Check truth table compliance
-- - Validate timing constraints and requirements
-- - Prove functional equivalence between architectures
--
-- ASSERTION-BASED VERIFICATION:
-- - Assert correct selection behavior
-- - Check for proper output assignment
-- - Verify no undefined output states
-- - Validate timing relationships
-- - Check select signal decode correctness
--
-- ============================================================================
-- COMPARISON WITH OTHER MULTIPLEXERS:
-- ============================================================================
--
-- 2-TO-1 vs 4-TO-1 MULTIPLEXER:
-- - 2-to-1: 1 select bit, simpler logic
-- - 4-to-1: 2 select bits, more complex decode
-- - 4-to-1 more versatile for multiple options
-- - 2-to-1 more efficient for binary selection
--
-- RESOURCE COMPARISON:
-- - 4-to-1 MUX: 1 LUT in modern FPGAs
-- - 8-to-1 MUX: 2 LUTs (or 1 LUT7/8)
-- - 16-to-1 MUX: Multiple LUTs, tree structure
-- - Choice depends on application requirements
--
-- PERFORMANCE COMPARISON:
-- - 4-to-1 MUX: Minimal propagation delay
-- - Larger MUX: Logarithmic delay increase
-- - Tree structure affects timing
-- - Consider critical path requirements
--
-- COMPLEXITY COMPARISON:
-- - 4-to-1: Moderate complexity, good balance
-- - 2-to-1: Simple but limited functionality
-- - 8-to-1+: Higher complexity, more versatile
-- - Sweet spot for many applications
--
-- ============================================================================
-- MULTIPLEXER DESIGN PATTERNS:
-- ============================================================================
--
-- BASIC SELECTION PATTERN:
-- - Simple input selection based on control
-- - Most common multiplexer usage
-- - Direct implementation of selection logic
-- - Suitable for most applications
--
-- HIERARCHICAL PATTERN:
-- - Build from smaller multiplexers
-- - Modular and scalable design
-- - Easy to understand and maintain
-- - Good for complex routing requirements
--
-- PARAMETERIZED PATTERN:
-- - Generic multiplexer with configurable inputs
-- - Use generics for input count and width
-- - Reusable component design
-- - Suitable for library development
--
-- PIPELINE PATTERN:
-- - Add registers for high-speed operation
-- - Break critical paths with flip-flops
-- - Increase throughput at cost of latency
-- - Suitable for high-frequency designs
--
-- PRIORITY PATTERN:
-- - Implement priority-based selection
-- - Handle multiple active inputs
-- - Add conflict resolution logic
-- - Suitable for interrupt controllers
--
-- ============================================================================
-- IMPLEMENTATION TEMPLATE:
-- ============================================================================
--
-- [Add your library declarations here]
--
-- [Add your entity declaration here]
--
-- [Add your architecture implementation here]
--
-- ============================================================================