-- ============================================================================
-- Up/Down Counter Implementation - Programming Guidance
-- ============================================================================
-- 
-- PROJECT OVERVIEW:
-- This file implements an up/down counter, a versatile sequential circuit that
-- can count in both ascending and descending directions based on a control
-- signal. Up/down counters are essential components in digital systems for
-- bidirectional counting, position tracking, and control applications.
--
-- LEARNING OBJECTIVES:
-- 1. Understand bidirectional counting principles
-- 2. Learn control signal implementation for direction
-- 3. Practice parameterized counter design
-- 4. Explore overflow/underflow handling
-- 5. Understand applications in control systems
--
-- ============================================================================
-- STEP-BY-STEP IMPLEMENTATION GUIDE:
-- ============================================================================
--
-- STEP 1: LIBRARY DECLARATIONS
-- ----------------------------------------------------------------------------
-- Required Libraries:
-- - IEEE library for standard logic types
-- - std_logic_1164 package for std_logic and std_logic_vector
-- - numeric_std package for arithmetic operations
-- 
-- TODO: Add library IEEE;
-- TODO: Add use IEEE.std_logic_1164.all;
-- TODO: Add use IEEE.numeric_std.all;
--
-- ============================================================================
-- STEP 2: ENTITY DECLARATION
-- ============================================================================
-- The entity defines the interface for the up/down counter
--
-- Entity Requirements:
-- - Name: up_down_counter (maintain current naming convention)
-- - Generic parameters for width and modulus
-- - Inputs: clock, reset, enable, up_down, load, data
-- - Outputs: count, overflow, underflow, terminal_count
--
-- Generic Parameters:
-- - WIDTH : positive := 4 (Counter bit width)
-- - MAX_COUNT : positive := 15 (Maximum count value)
-- - MIN_COUNT : natural := 0 (Minimum count value)
--
-- Port Specifications:
-- - clk : in std_logic (Clock input for synchronous operation)
-- - reset : in std_logic (Reset signal - active high)
-- - enable : in std_logic (Enable signal for counting)
-- - up_down : in std_logic (Direction control: '1' = up, '0' = down)
-- - load : in std_logic (Load control for parallel loading)
-- - load_data : in std_logic_vector(WIDTH-1 downto 0) (Parallel load data)
-- - count : out std_logic_vector(WIDTH-1 downto 0) (Current count value)
-- - overflow : out std_logic (Overflow flag - count exceeded maximum)
-- - underflow : out std_logic (Underflow flag - count below minimum)
-- - terminal_count : out std_logic (Terminal count reached)
--
-- Optional Ports:
-- - carry_in : in std_logic (Carry input for cascading)
-- - carry_out : out std_logic (Carry output for cascading)
-- - borrow_in : in std_logic (Borrow input for cascading)
-- - borrow_out : out std_logic (Borrow output for cascading)
-- - preset : in std_logic (Preset signal - active high)
-- - clear : in std_logic (Clear signal - active high)
--
-- Design Considerations:
-- - Parameterizable width and range
-- - Bidirectional counting capability
-- - Overflow/underflow detection
-- - Parallel load functionality
-- - Cascading support
-- - Control signal priorities
--
-- TODO: Declare entity with appropriate generics and ports
-- TODO: Add comprehensive port comments
-- TODO: Consider optional features needed
-- TODO: Plan for cascading requirements
--
-- ============================================================================
-- STEP 3: UP/DOWN COUNTER OPERATION DEFINITIONS
-- ============================================================================
--
-- UP/DOWN COUNTER PRINCIPLES:
-- - Count up when up_down = '1'
-- - Count down when up_down = '0'
-- - Enable control for conditional counting
-- - Parallel load capability
-- - Overflow/underflow detection
-- - Modular arithmetic operation
--
-- OPERATION TABLE (Basic Up/Down Counter):
-- Clock | Reset | Enable | Up_Down | Load | Operation
-- ------|-------|--------|---------|------|----------
--   X   |   1   |   X    |    X    |  X   | Reset to MIN_COUNT
--   ↑   |   0   |   0    |    X    |  X   | Hold current count
--   ↑   |   0   |   1    |    X    |  1   | Load parallel data
--   ↑   |   0   |   1    |    1    |  0   | Count up
--   ↑   |   0   |   1    |    0    |  0   | Count down
--
-- COUNTING BEHAVIOR:
-- - Up counting: count <= count + 1 (with overflow check)
-- - Down counting: count <= count - 1 (with underflow check)
-- - Modular operation: wrap around at boundaries
-- - Load operation: count <= load_data
-- - Reset operation: count <= MIN_COUNT
--
-- OVERFLOW/UNDERFLOW CONDITIONS:
-- - Overflow: count = MAX_COUNT and up_down = '1' and enable = '1'
-- - Underflow: count = MIN_COUNT and up_down = '0' and enable = '1'
-- - Wrap-around behavior on overflow/underflow
-- - Flag generation for external monitoring
--
-- TERMINAL COUNT CONDITIONS:
-- - Up counting: terminal_count when count = MAX_COUNT
-- - Down counting: terminal_count when count = MIN_COUNT
-- - Used for cascading multiple counters
-- - Enables higher-order counter stages
--
-- TIMING REQUIREMENTS:
-- - Setup time: Control signals stable before clock edge
-- - Hold time: Control signals stable after clock edge
-- - Clock-to-Q delay: Time from clock to output change
-- - Reset recovery time: Time from reset release to clock
-- - Load data setup time: Data stable before load
--
-- TODO: Define operation tables for chosen configuration
-- TODO: Specify overflow/underflow behavior
-- TODO: Plan terminal count generation
-- TODO: Consider cascading requirements
--
-- ============================================================================
-- STEP 4: ARCHITECTURE IMPLEMENTATION OPTIONS
-- ============================================================================
--
-- OPTION 1: BASIC SYNCHRONOUS UP/DOWN COUNTER
-- ----------------------------------------------------------------------------
-- Simple up/down counter with basic functionality
--
-- Implementation Approach:
-- - Single process for synchronous operation
-- - Conditional increment/decrement logic
-- - Synchronous reset functionality
-- - Basic overflow/underflow detection
--
-- Example Structure:
-- architecture behavioral of up_down_counter is
--     signal count_internal : unsigned(WIDTH-1 downto 0) := (others => '0');
--     signal overflow_internal : std_logic := '0';
--     signal underflow_internal : std_logic := '0';
-- begin
--     -- Up/Down counter process
--     counter_proc: process(clk)
--     begin
--         if rising_edge(clk) then
--             if reset = '1' then
--                 count_internal <= to_unsigned(MIN_COUNT, WIDTH);
--                 overflow_internal <= '0';
--                 underflow_internal <= '0';
--             elsif enable = '1' then
--                 if up_down = '1' then
--                     -- Count up
--                     if count_internal = MAX_COUNT then
--                         count_internal <= to_unsigned(MIN_COUNT, WIDTH);
--                         overflow_internal <= '1';
--                     else
--                         count_internal <= count_internal + 1;
--                         overflow_internal <= '0';
--                     end if;
--                     underflow_internal <= '0';
--                 else
--                     -- Count down
--                     if count_internal = MIN_COUNT then
--                         count_internal <= to_unsigned(MAX_COUNT, WIDTH);
--                         underflow_internal <= '1';
--                     else
--                         count_internal <= count_internal - 1;
--                         underflow_internal <= '0';
--                     end if;
--                     overflow_internal <= '0';
--                 end if;
--             end if;
--         end if;
--     end process;
--     
--     -- Output assignments
--     count <= std_logic_vector(count_internal);
--     overflow <= overflow_internal;
--     underflow <= underflow_internal;
--     terminal_count <= '1' when (count_internal = MAX_COUNT and up_down = '1') or
--                               (count_internal = MIN_COUNT and up_down = '0') else '0';
-- end behavioral;
--
-- Counting Logic Explanation:
-- - Up counting: increment with overflow check
-- - Down counting: decrement with underflow check
-- - Wrap-around behavior at boundaries
-- - Flag generation for monitoring
--
-- Advantages:
-- - Simple implementation
-- - Predictable behavior
-- - Low resource usage
-- - Easy to understand
--
-- Disadvantages:
-- - No parallel load capability
-- - No asynchronous reset
-- - Limited control features
-- - No cascading support
--
-- TODO: Implement basic up/down counter
-- TODO: Verify counting directions
-- TODO: Test overflow/underflow behavior
-- TODO: Validate terminal count generation
--
-- OPTION 2: FULL-FEATURED UP/DOWN COUNTER
-- ----------------------------------------------------------------------------
-- Comprehensive up/down counter with all features
--
-- Implementation Approach:
-- - Parallel load capability
-- - Asynchronous reset option
-- - Comprehensive flag generation
-- - Cascading support
--
-- Example Structure:
-- architecture full_featured of up_down_counter is
--     signal count_internal : unsigned(WIDTH-1 downto 0) := to_unsigned(MIN_COUNT, WIDTH);
--     signal overflow_internal : std_logic := '0';
--     signal underflow_internal : std_logic := '0';
--     signal terminal_count_internal : std_logic := '0';
-- begin
--     -- Full-featured up/down counter process
--     counter_proc: process(clk, reset)
--     begin
--         if reset = '1' then
--             count_internal <= to_unsigned(MIN_COUNT, WIDTH);
--             overflow_internal <= '0';
--             underflow_internal <= '0';
--         elsif rising_edge(clk) then
--             -- Clear flags by default
--             overflow_internal <= '0';
--             underflow_internal <= '0';
--             
--             if load = '1' then
--                 -- Parallel load operation
--                 count_internal <= unsigned(load_data);
--             elsif enable = '1' then
--                 if up_down = '1' then
--                     -- Count up with carry
--                     if count_internal = MAX_COUNT then
--                         count_internal <= to_unsigned(MIN_COUNT, WIDTH);
--                         overflow_internal <= '1';
--                     else
--                         count_internal <= count_internal + 1;
--                     end if;
--                 else
--                     -- Count down with borrow
--                     if count_internal = MIN_COUNT then
--                         count_internal <= to_unsigned(MAX_COUNT, WIDTH);
--                         underflow_internal <= '1';
--                     else
--                         count_internal <= count_internal - 1;
--                     end if;
--                 end if;
--             end if;
--         end if;
--     end process;
--     
--     -- Terminal count generation
--     terminal_count_internal <= '1' when (count_internal = MAX_COUNT and up_down = '1') or
--                                        (count_internal = MIN_COUNT and up_down = '0') else '0';
--     
--     -- Output assignments
--     count <= std_logic_vector(count_internal);
--     overflow <= overflow_internal;
--     underflow <= underflow_internal;
--     terminal_count <= terminal_count_internal;
-- end full_featured;
--
-- Control Signal Priority (highest to lowest):
-- 1. Asynchronous Reset (forces count to MIN_COUNT)
-- 2. Parallel Load (loads external data)
-- 3. Count Enable (allows counting operation)
-- 4. Hold current count (default)
--
-- Parallel Load Features:
-- - Immediate data loading
-- - Overrides counting operation
-- - Useful for initialization
-- - Supports preset values
--
-- Advantages:
-- - Complete functionality
-- - Professional features
-- - Flexible operation modes
-- - Industry-standard interface
--
-- Disadvantages:
-- - Complex control logic
-- - Higher resource usage
-- - More complex verification
-- - Potential timing issues
--
-- TODO: Implement full-featured up/down counter
-- TODO: Add parallel load functionality
-- TODO: Test all control combinations
-- TODO: Verify flag generation
--
-- OPTION 3: CASCADABLE UP/DOWN COUNTER
-- ----------------------------------------------------------------------------
-- Up/down counter designed for multi-stage cascading
--
-- Implementation Approach:
-- - Carry/borrow chain support
-- - Ripple or synchronous cascading
-- - Terminal count propagation
-- - Multi-stage coordination
--
-- Example Structure:
-- architecture cascadable of up_down_counter is
--     signal count_internal : unsigned(WIDTH-1 downto 0) := to_unsigned(MIN_COUNT, WIDTH);
--     signal carry_out_internal : std_logic := '0';
--     signal borrow_out_internal : std_logic := '0';
--     signal enable_internal : std_logic;
-- begin
--     -- Enable logic for cascading
--     enable_internal <= enable and ((carry_in and up_down) or (borrow_in and not up_down));
--     
--     -- Cascadable up/down counter process
--     counter_proc: process(clk, reset)
--     begin
--         if reset = '1' then
--             count_internal <= to_unsigned(MIN_COUNT, WIDTH);
--             carry_out_internal <= '0';
--             borrow_out_internal <= '0';
--         elsif rising_edge(clk) then
--             -- Clear carry/borrow by default
--             carry_out_internal <= '0';
--             borrow_out_internal <= '0';
--             
--             if load = '1' then
--                 count_internal <= unsigned(load_data);
--             elsif enable_internal = '1' then
--                 if up_down = '1' then
--                     -- Count up with carry generation
--                     if count_internal = MAX_COUNT then
--                         count_internal <= to_unsigned(MIN_COUNT, WIDTH);
--                         carry_out_internal <= '1';
--                     else
--                         count_internal <= count_internal + 1;
--                     end if;
--                 else
--                     -- Count down with borrow generation
--                     if count_internal = MIN_COUNT then
--                         count_internal <= to_unsigned(MAX_COUNT, WIDTH);
--                         borrow_out_internal <= '1';
--                     else
--                         count_internal <= count_internal - 1;
--                     end if;
--                 end if;
--             end if;
--         end if;
--     end process;
--     
--     -- Output assignments
--     count <= std_logic_vector(count_internal);
--     carry_out <= carry_out_internal;
--     borrow_out <= borrow_out_internal;
--     terminal_count <= '1' when (count_internal = MAX_COUNT and up_down = '1') or
--                               (count_internal = MIN_COUNT and up_down = '0') else '0';
-- end cascadable;
--
-- Cascading Features:
-- - Carry/borrow chain propagation
-- - Multi-stage counter support
-- - Ripple or synchronous operation
-- - Scalable bit width
--
-- Carry/Borrow Logic:
-- - Carry out: generated on overflow during up counting
-- - Borrow out: generated on underflow during down counting
-- - Carry/borrow in: enables counting from previous stage
-- - Chain coordination for large counters
--
-- Advantages:
-- - Scalable architecture
-- - Multi-stage support
-- - Flexible bit width
-- - Standard cascading interface
--
-- Disadvantages:
-- - Complex cascading logic
-- - Timing considerations
-- - Propagation delays
-- - Design complexity
--
-- TODO: Implement cascadable up/down counter
-- TODO: Add carry/borrow logic
-- TODO: Test cascading operation
-- TODO: Verify multi-stage behavior
--
-- OPTION 4: PARAMETERIZED MODULAR COUNTER
-- ----------------------------------------------------------------------------
-- Highly parameterized counter with configurable modulus
--
-- Implementation Approach:
-- - Generic parameters for full customization
-- - Configurable count range
-- - Modular arithmetic
-- - Flexible boundary conditions
--
-- Example Structure:
-- architecture parameterized of up_down_counter is
--     constant COUNT_RANGE : positive := MAX_COUNT - MIN_COUNT + 1;
--     signal count_internal : unsigned(WIDTH-1 downto 0) := to_unsigned(MIN_COUNT, WIDTH);
--     signal next_count : unsigned(WIDTH-1 downto 0);
-- begin
--     -- Next count calculation
--     next_count_proc: process(count_internal, up_down, enable)
--     begin
--         if enable = '1' then
--             if up_down = '1' then
--                 -- Up counting with modular arithmetic
--                 if count_internal = MAX_COUNT then
--                     next_count <= to_unsigned(MIN_COUNT, WIDTH);
--                 else
--                     next_count <= count_internal + 1;
--                 end if;
--             else
--                 -- Down counting with modular arithmetic
--                 if count_internal = MIN_COUNT then
--                     next_count <= to_unsigned(MAX_COUNT, WIDTH);
--                 else
--                     next_count <= count_internal - 1;
--                 end if;
--             end if;
--         else
--             next_count <= count_internal;
--         end if;
--     end process;
--     
--     -- Counter register
--     counter_reg: process(clk, reset)
--     begin
--         if reset = '1' then
--             count_internal <= to_unsigned(MIN_COUNT, WIDTH);
--         elsif rising_edge(clk) then
--             if load = '1' then
--                 count_internal <= unsigned(load_data);
--             else
--                 count_internal <= next_count;
--             end if;
--         end if;
--     end process;
--     
--     -- Flag generation
--     overflow <= '1' when (count_internal = MAX_COUNT and up_down = '1' and enable = '1') else '0';
--     underflow <= '1' when (count_internal = MIN_COUNT and up_down = '0' and enable = '1') else '0';
--     terminal_count <= '1' when (count_internal = MAX_COUNT and up_down = '1') or
--                               (count_internal = MIN_COUNT and up_down = '0') else '0';
--     
--     -- Output assignment
--     count <= std_logic_vector(count_internal);
-- end parameterized;
--
-- Parameterization Benefits:
-- - Configurable count range
-- - Flexible modulus selection
-- - Reusable component
-- - Technology independent
--
-- Modular Arithmetic:
-- - Wrap-around at boundaries
-- - Configurable range limits
-- - Efficient implementation
-- - Predictable behavior
--
-- Advantages:
-- - Highly configurable
-- - Reusable design
-- - Efficient implementation
-- - Clear separation of concerns
--
-- Disadvantages:
-- - Complex parameterization
-- - Generic validation needed
-- - Synthesis considerations
-- - Documentation requirements
--
-- TODO: Implement parameterized counter
-- TODO: Validate generic parameters
-- TODO: Test modular arithmetic
-- TODO: Verify configurability
--
-- ============================================================================
-- STEP 5: ADVANCED UP/DOWN COUNTER FEATURES
-- ============================================================================
--
-- GRAY CODE COUNTING:
-- - Non-binary counting sequence
-- - Single bit change per transition
-- - Reduced switching noise
-- - Asynchronous interface compatibility
--
-- JOHNSON COUNTER INTEGRATION:
-- - Ring counter with feedback
-- - Self-decoding outputs
-- - Reduced decode logic
-- - Specific sequence generation
--
-- PRESCALER FUNCTIONALITY:
-- - Programmable division ratios
-- - Clock frequency reduction
-- - Timing reference generation
-- - System clock management
--
-- BCD COUNTING MODE:
-- - Binary-coded decimal operation
-- - Decimal display compatibility
-- - Modulo-10 operation
-- - Human-readable output
--
-- TODO: Select appropriate advanced features
-- TODO: Implement chosen enhancements
-- TODO: Verify advanced functionality
-- TODO: Test integration capabilities
--
-- ============================================================================
-- IMPLEMENTATION CONSIDERATIONS:
-- ============================================================================
--
-- GENERIC PARAMETER VALIDATION:
-- - Width range checking
-- - Count range validation
-- - Consistency verification
-- - Error handling
--
-- ARITHMETIC OVERFLOW HANDLING:
-- - Boundary condition management
-- - Wrap-around behavior
-- - Flag generation timing
-- - Cascading implications
--
-- TIMING OPTIMIZATION:
-- - Critical path analysis
-- - Pipeline considerations
-- - Clock frequency optimization
-- - Setup/hold margin
--
-- SYNTHESIS OPTIMIZATION:
-- - Resource utilization
-- - Timing constraints
-- - Power optimization
-- - Area minimization
--
-- TESTABILITY:
-- - Scan chain integration
-- - Test pattern generation
-- - Fault coverage analysis
-- - Built-in self-test
--
-- ============================================================================
-- APPLICATIONS:
-- ============================================================================
--
-- 1. POSITION CONTROL:
--    - Motor position tracking
--    - Encoder interface
--    - Bidirectional movement
--    - Position feedback
--
-- 2. DIGITAL FILTERS:
--    - Address generation
--    - Delay line control
--    - Sample indexing
--    - Buffer management
--
-- 3. COMMUNICATION PROTOCOLS:
--    - Frame counting
--    - Sequence numbering
--    - Error detection
--    - Flow control
--
-- 4. MEMORY INTERFACES:
--    - Address generation
--    - Bank switching
--    - Refresh counting
--    - Access control
--
-- 5. CONTROL SYSTEMS:
--    - State sequencing
--    - Event counting
--    - Timing control
--    - Process monitoring
--
-- ============================================================================
-- TESTING STRATEGY:
-- ============================================================================
--
-- FUNCTIONAL TESTING:
-- - Verify up counting operation
-- - Test down counting operation
-- - Check direction control
-- - Validate enable functionality
-- - Test parallel load operation
-- - Verify reset behavior
--
-- BOUNDARY TESTING:
-- - Test overflow conditions
-- - Verify underflow behavior
-- - Check wrap-around operation
-- - Validate terminal count generation
-- - Test boundary transitions
--
-- CONTROL SIGNAL TESTING:
-- - Test all control combinations
-- - Verify signal priorities
-- - Check simultaneous assertions
-- - Validate timing relationships
-- - Test edge cases
--
-- CASCADING TESTING:
-- - Multi-stage operation
-- - Carry/borrow propagation
-- - Synchronization verification
-- - Performance analysis
-- - Scalability testing
--
-- STRESS TESTING:
-- - Continuous operation
-- - High-frequency counting
-- - Temperature variation
-- - Voltage variation
-- - Long-term reliability
--
-- ============================================================================
-- RECOMMENDED IMPLEMENTATION APPROACH:
-- ============================================================================
--
-- FOR BEGINNERS:
-- 1. Start with basic up/down counter
-- 2. Implement direction control
-- 3. Add enable functionality
-- 4. Test counting operations
-- 5. Verify overflow/underflow
--
-- FOR INTERMEDIATE USERS:
-- 1. Add parallel load capability
-- 2. Implement flag generation
-- 3. Create comprehensive testbench
-- 4. Optimize for target technology
-- 5. Add cascading support
--
-- FOR ADVANCED USERS:
-- 1. Implement parameterized version
-- 2. Add advanced features
-- 3. Create library-quality component
-- 4. Implement power optimizations
-- 5. Develop production verification suite
--
-- ============================================================================
-- EXTENSION EXERCISES:
-- ============================================================================
--
-- 1. MULTI-STAGE COUNTER:
--    - Chain multiple counters
--    - Synchronous operation
--    - Carry/borrow propagation
--    - Large bit width support
--
-- 2. PROGRAMMABLE COUNTER:
--    - Runtime modulus configuration
--    - Dynamic range adjustment
--    - Control register interface
--    - Flexible operation modes
--
-- 3. GRAY CODE COUNTER:
--    - Non-binary sequence
--    - Single bit transitions
--    - Asynchronous compatibility
--    - Noise reduction
--
-- 4. BCD UP/DOWN COUNTER:
--    - Decimal counting
--    - Display compatibility
--    - Modulo-10 operation
--    - Multi-digit support
--
-- 5. FREQUENCY SYNTHESIZER:
--    - Programmable division
--    - Fractional ratios
--    - Phase accumulation
--    - Clock generation
--
-- ============================================================================
-- COMMON MISTAKES TO AVOID:
-- ============================================================================
--
-- 1. BOUNDARY CONDITION ERRORS:
--    - Incorrect overflow detection
--    - Wrong underflow handling
--    - Boundary value mistakes
--    - Wrap-around errors
--
-- 2. CONTROL SIGNAL CONFLICTS:
--    - Priority resolution issues
--    - Simultaneous assertion problems
--    - Timing relationship errors
--    - Enable logic mistakes
--
-- 3. ARITHMETIC IMPLEMENTATION ERRORS:
--    - Type conversion mistakes
--    - Range checking oversights
--    - Modular arithmetic errors
--    - Carry/borrow logic flaws
--
-- 4. PARAMETERIZATION ISSUES:
--    - Generic validation missing
--    - Range checking inadequate
--    - Consistency verification lacking
--    - Default value problems
--
-- 5. SYNTHESIS OPTIMIZATION OVERSIGHTS:
--    - Resource utilization inefficiency
--    - Timing constraint violations
--    - Power optimization missed
--    - Technology mapping issues
--
-- ============================================================================
-- DESIGN VERIFICATION CHECKLIST:
-- ============================================================================
--
-- □ Entity declaration with proper generics and ports
-- □ Up counting operation working correctly
-- □ Down counting operation functioning properly
-- □ Direction control working as expected
-- □ Enable functionality implemented correctly
-- □ Parallel load operation verified
-- □ Reset functionality working properly
-- □ Overflow detection accurate
-- □ Underflow detection correct
-- □ Terminal count generation proper
-- □ Wrap-around behavior correct
-- □ Control signal priorities right
-- □ Cascading support functional (if implemented)
-- □ Flag generation timing correct
-- □ Generic parameter validation complete
-- □ Synthesis results acceptable
-- □ Resource utilization optimized
-- □ Testbench covers all scenarios
-- □ Edge cases thoroughly tested
-- □ Documentation complete and accurate
-- □ Code follows design standards
-- □ Performance requirements met
--
-- ============================================================================
-- DIGITAL DESIGN CONTEXT:
-- ============================================================================
--
-- RELATIONSHIP TO OTHER COUNTERS:
-- - Binary Counter: Subset with fixed direction
-- - Ring Counter: Different counting sequence
-- - Johnson Counter: Modified ring counter
-- - Gray Counter: Non-binary sequence
--
-- SEQUENTIAL LOGIC PRINCIPLES:
-- - State-based operation
-- - Clock synchronization
-- - Memory element behavior
-- - Timing relationships
--
-- SYSTEM INTEGRATION ASPECTS:
-- - Control system design
-- - Position tracking systems
-- - Communication protocols
-- - Memory management
--
-- ============================================================================
-- PHYSICAL IMPLEMENTATION NOTES:
-- ============================================================================
--
-- FPGA IMPLEMENTATION:
-- - Efficient counter utilization
-- - Clock network optimization
-- - Reset distribution
-- - Timing constraint application
--
-- ASIC IMPLEMENTATION:
-- - Standard cell selection
-- - Custom cell opportunities
-- - Layout optimization
-- - Power grid considerations
--
-- PERFORMANCE CHARACTERISTICS:
-- - Frequency scaling behavior
-- - Power consumption patterns
-- - Area utilization
-- - Temperature sensitivity
--
-- ============================================================================
-- ADVANCED CONCEPTS:
-- ============================================================================
--
-- MODULAR ARITHMETIC:
-- - Wrap-around behavior
-- - Boundary conditions
-- - Range validation
-- - Efficiency optimization
--
-- CASCADING TECHNIQUES:
-- - Ripple vs synchronous
-- - Carry/borrow chains
-- - Multi-stage coordination
-- - Timing considerations
--
-- POWER MANAGEMENT:
-- - Clock gating strategies
-- - Activity-based optimization
-- - Dynamic power scaling
-- - Leakage reduction
--
-- ============================================================================
-- SIMULATION AND VERIFICATION NOTES:
-- ============================================================================
--
-- TESTBENCH DEVELOPMENT:
-- - Comprehensive test scenarios
-- - Automated verification
-- - Coverage analysis
-- - Performance measurement
--
-- VERIFICATION METHODOLOGY:
-- - Functional verification
-- - Timing verification
-- - Power verification
-- - Reliability verification
--
-- DEBUGGING TECHNIQUES:
-- - Waveform analysis
-- - State transition tracing
-- - Timing analysis
-- - Resource utilization analysis
--
-- ============================================================================
-- IMPLEMENTATION TEMPLATE:
-- ============================================================================
--
-- [Add your library declarations here]
--
-- [Add your entity declaration here with generics]
--
-- [Add your architecture implementation here]
--
-- ============================================================================