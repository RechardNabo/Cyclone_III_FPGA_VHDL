-- ============================================================================
-- PCI Bridge FSMD (FSM + Datapath) - Programming Guidance
-- ============================================================================
--
-- PROJECT OVERVIEW:
-- This header documents an integrated FSMD design for a PCI(-like) bridge.
-- State actions explicitly drive datapath transfers (registers/FIFOs/muxes),
-- producing a single, coherent implementation while maintaining clean signal
-- partitioning.
--
-- LEARNING OBJECTIVES:
-- - Map protocol phases to state-driven register/FIFO operations
-- - Keep datapath enables and mux selects derived from states
-- - Maintain testability with clear defaults and handshakes
--
-- IMPLEMENTATION GUIDE:
-- 1) LIBRARIES
--    TODO: library IEEE;
--    TODO: use IEEE.std_logic_1164.all;
--    TODO: use IEEE.numeric_std.all;
--
-- 2) ENTITY (FSMD INTERFACE)
--    Typical ports:
--    - clk, reset : in std_logic
--    - start, rw  : in std_logic
--    - addr_in    : in unsigned(ADDR_WIDTH-1 downto 0)
--    - wdata_in   : in unsigned(DATA_WIDTH-1 downto 0)
--    - rdata_out  : out unsigned(DATA_WIDTH-1 downto 0)
--    - empty, full, ready : in std_logic
--    - push, pop, drive_en : out std_logic
--    - done, error : out std_logic
--    Generics: ADDR_WIDTH := 32, DATA_WIDTH := 32
--
-- 3) STATE/ACTION EXAMPLE
--    - IDLE: defaults, clear enables
--    - ADDRESS: latch addr_in
--    - DATA_WR: push wdata_in to write FIFO
--    - DATA_RD: pop from read FIFO → rdata_out
--    - COMPLETE: assert done
--
-- 4) CODING STYLE
--    - Single clocked state register
--    - Combinational next-state + control generation
--    - Datapath transfers gated by current state
--    - Defaults provided to avoid inferred latches
--
-- 5) TESTING
--    - FIFO underflow/overflow protection
--    - Latency counters and ready behavior
--    - Back-to-back transaction coverage
--
-- Use this header as a blueprint for the integrated architecture, then add
-- detailed signals, counters, and handshakes per your protocol.
-- ============================================================================