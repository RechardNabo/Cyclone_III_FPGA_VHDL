-- ============================================================================
-- Priority Encoder Implementation - Programming Guidance
-- ============================================================================
-- 
-- PROJECT OVERVIEW:
-- This file implements a priority encoder, a combinational circuit that encodes
-- the position of the highest priority active input into a binary code. Priority
-- encoders are essential components in interrupt controllers, arbitration circuits,
-- and resource allocation systems. They provide a systematic way to handle
-- multiple simultaneous requests by establishing a priority hierarchy.
--
-- LEARNING OBJECTIVES:
-- 1. Understand priority encoding principles and applications
-- 2. Learn binary encoding techniques for position representation
-- 3. Practice hierarchical priority resolution logic
-- 4. Explore cascading methods for larger input sets
-- 5. Understand interrupt controller and arbitration applications
--
-- ============================================================================
-- STEP-BY-STEP IMPLEMENTATION GUIDE:
-- ============================================================================
--
-- STEP 1: LIBRARY DECLARATIONS
-- ----------------------------------------------------------------------------
-- Required Libraries:
-- - IEEE library for standard logic types
-- - std_logic_1164 package for std_logic and logical operators
-- - numeric_std package for arithmetic operations (recommended)
-- - std_logic_arith and std_logic_unsigned (alternative, not recommended)
-- 
-- TODO: Add library IEEE;
-- TODO: Add use IEEE.std_logic_1164.all;
-- TODO: Add use IEEE.numeric_std.all; (recommended approach)
-- TODO: Consider use IEEE.std_logic_arith.all; (alternative approach)
--
-- ============================================================================
-- STEP 2: ENTITY DECLARATION
-- ============================================================================
-- The entity defines the interface for the priority encoder
--
-- Entity Requirements:
-- - Name: priority_encoder (maintain current naming convention)
-- - Inputs: Multiple request inputs, enable control
-- - Outputs: Encoded priority position, valid output flag
-- - Consider expandable design for different input counts
--
-- Port Specifications:
-- - Requests : in std_logic_vector(7 downto 0) (Input requests - 8 inputs)
-- - Enable : in std_logic (Encoder enable signal)
-- - Encoded_Output : out std_logic_vector(2 downto 0) (3-bit encoded position)
-- - Valid_Output : out std_logic (Valid encoding flag)
-- - Any_Request : out std_logic (Any input active flag - optional)
--
-- Priority Convention:
-- - Higher index = Higher priority (Request(7) has highest priority)
-- - Lower index = Lower priority (Request(0) has lowest priority)
-- - Alternative: Lower index = Higher priority (design choice)
--
-- TODO: Declare entity with appropriate port names
-- TODO: Add detailed port comments
-- TODO: Consider signal naming conventions
-- TODO: Plan for different input counts (16, 32, 64 inputs)
--
-- ============================================================================
-- STEP 3: PRIORITY ENCODING OPERATION DEFINITIONS
-- ============================================================================
--
-- PRIORITY ENCODING PRINCIPLE:
-- - Scan inputs from highest to lowest priority
-- - Encode position of first (highest priority) active input
-- - Ignore all lower priority active inputs
-- - Generate valid flag when any input is active
--
-- ENCODING TABLE (8-input example, MSB has highest priority):
-- Requests[7:0] | Encoded_Output[2:0] | Valid_Output | Priority Input
-- 1xxxxxxx      | 111                 | 1            | Request(7)
-- 01xxxxxx      | 110                 | 1            | Request(6)
-- 001xxxxx      | 101                 | 1            | Request(5)
-- 0001xxxx      | 100                 | 1            | Request(4)
-- 00001xxx      | 011                 | 1            | Request(3)
-- 000001xx      | 010                 | 1            | Request(2)
-- 0000001x      | 001                 | 1            | Request(1)
-- 00000001      | 000                 | 1            | Request(0)
-- 00000000      | XXX                 | 0            | No request
--
-- ALTERNATIVE ENCODING (LSB has highest priority):
-- Requests[7:0] | Encoded_Output[2:0] | Valid_Output | Priority Input
-- xxxxxxx1      | 000                 | 1            | Request(0)
-- xxxxxx10      | 001                 | 1            | Request(1)
-- xxxxx100      | 010                 | 1            | Request(2)
-- xxxx1000      | 011                 | 1            | Request(3)
-- xxx10000      | 100                 | 1            | Request(4)
-- xx100000      | 101                 | 1            | Request(5)
-- x1000000      | 110                 | 1            | Request(6)
-- 10000000      | 111                 | 1            | Request(7)
-- 00000000      | XXX                 | 0            | No request
--
-- OUTPUT CHARACTERISTICS:
-- - Encoded_Output: Binary representation of highest priority active input
-- - Valid_Output: '1' when at least one input is active, '0' otherwise
-- - Any_Request: Optional output indicating any request present
--
-- TODO: Define priority encoding truth table
-- TODO: Document priority convention choice
-- TODO: Plan for output encoding format
-- TODO: Consider don't-care optimization opportunities
--
-- ============================================================================
-- STEP 4: ARCHITECTURE IMPLEMENTATION OPTIONS
-- ============================================================================
--
-- OPTION 1: BEHAVIORAL ARCHITECTURE (IF-THEN-ELSE CASCADE)
-- ----------------------------------------------------------------------------
-- Use priority-ordered conditional statements
--
-- Implementation Approach:
-- - Use process with if-then-elsif cascade
-- - Check inputs from highest to lowest priority
-- - First active input determines output
-- - Simple and readable implementation
--
-- Example Structure (MSB highest priority):
-- process(Requests, Enable)
-- begin
--     if Enable = '1' then
--         if Requests(7) = '1' then
--             Encoded_Output <= "111";
--             Valid_Output <= '1';
--         elsif Requests(6) = '1' then
--             Encoded_Output <= "110";
--             Valid_Output <= '1';
--         elsif Requests(5) = '1' then
--             Encoded_Output <= "101";
--             Valid_Output <= '1';
--         elsif Requests(4) = '1' then
--             Encoded_Output <= "100";
--             Valid_Output <= '1';
--         elsif Requests(3) = '1' then
--             Encoded_Output <= "011";
--             Valid_Output <= '1';
--         elsif Requests(2) = '1' then
--             Encoded_Output <= "010";
--             Valid_Output <= '1';
--         elsif Requests(1) = '1' then
--             Encoded_Output <= "001";
--             Valid_Output <= '1';
--         elsif Requests(0) = '1' then
--             Encoded_Output <= "000";
--             Valid_Output <= '1';
--         else
--             Encoded_Output <= "000"; -- or don't care
--             Valid_Output <= '0';
--         end if;
--     else
--         Encoded_Output <= "000";
--         Valid_Output <= '0';
--     end if;
-- end process;
--
-- TODO: Implement behavioral architecture with if-then-elsif
-- TODO: Handle enable control logic
-- TODO: Verify priority ordering
-- TODO: Test synthesis results
--
-- OPTION 2: DATAFLOW ARCHITECTURE (CONCURRENT ASSIGNMENTS)
-- ----------------------------------------------------------------------------
-- Use concurrent signal assignments with conditional operators
--
-- Implementation Approach:
-- - Create intermediate priority signals
-- - Use conditional assignments for encoding
-- - Generate outputs concurrently
-- - Explicit logic for each condition
--
-- Example Structure:
-- -- Priority detection (MSB highest priority)
-- priority_7 <= Requests(7);
-- priority_6 <= Requests(6) and not Requests(7);
-- priority_5 <= Requests(5) and not (Requests(7) or Requests(6));
-- priority_4 <= Requests(4) and not (Requests(7) or Requests(6) or Requests(5));
-- priority_3 <= Requests(3) and not (Requests(7 downto 4) /= "0000");
-- priority_2 <= Requests(2) and not (Requests(7 downto 3) /= "00000");
-- priority_1 <= Requests(1) and not (Requests(7 downto 2) /= "000000");
-- priority_0 <= Requests(0) and not (Requests(7 downto 1) /= "0000000");
-- 
-- -- Encoding logic
-- Encoded_Output <= "111" when priority_7 = '1' else
--                   "110" when priority_6 = '1' else
--                   "101" when priority_5 = '1' else
--                   "100" when priority_4 = '1' else
--                   "011" when priority_3 = '1' else
--                   "010" when priority_2 = '1' else
--                   "001" when priority_1 = '1' else
--                   "000" when priority_0 = '1' else
--                   "000"; -- default case
-- 
-- Valid_Output <= (Requests /= "00000000") and Enable;
--
-- TODO: Implement dataflow architecture
-- TODO: Create priority detection signals
-- TODO: Implement concurrent encoding logic
-- TODO: Add enable gating
--
-- OPTION 3: STRUCTURAL ARCHITECTURE (HIERARCHICAL DESIGN)
-- ----------------------------------------------------------------------------
-- Use hierarchical components for scalable design
--
-- Implementation Approach:
-- - Create smaller priority encoder components
-- - Combine using tree structure
-- - Enable cascading for larger inputs
-- - Modular and scalable approach
--
-- Component Declarations:
-- component priority_encoder_4bit is
--     port (
--         Requests : in std_logic_vector(3 downto 0);
--         Enable : in std_logic;
--         Encoded_Output : out std_logic_vector(1 downto 0);
--         Valid_Output : out std_logic
--     );
-- end component;
--
-- Hierarchical Structure:
-- - Two 4-bit encoders for lower and upper halves
-- - Priority logic to select between halves
-- - Output multiplexing based on priority
-- - Additional bit for half selection
--
-- Signal Declarations:
-- signal lower_encoded, upper_encoded : std_logic_vector(1 downto 0);
-- signal lower_valid, upper_valid : std_logic;
-- signal upper_priority : std_logic;
--
-- TODO: Declare hierarchical components
-- TODO: Create tree structure for scalability
-- TODO: Implement output multiplexing
-- TODO: Handle cascading logic
--
-- OPTION 4: OPTIMIZED LOOP-BASED ARCHITECTURE
-- ----------------------------------------------------------------------------
-- Use for-loop for parameterized and compact implementation
--
-- Implementation Approach:
-- - Use for-loop to scan inputs
-- - Generate encoding using loop index
-- - Parameterizable for different input counts
-- - Compact and maintainable code
--
-- Example Structure:
-- process(Requests, Enable)
-- begin
--     Encoded_Output <= (others => '0');
--     Valid_Output <= '0';
--     
--     if Enable = '1' then
--         for i in Requests'high downto Requests'low loop
--             if Requests(i) = '1' then
--                 Encoded_Output <= std_logic_vector(to_unsigned(i, Encoded_Output'length));
--                 Valid_Output <= '1';
--                 exit; -- Exit on first (highest priority) match
--             end if;
--         end loop;
--     end if;
-- end process;
--
-- TODO: Implement loop-based architecture
-- TODO: Use generic parameters for scalability
-- TODO: Verify synthesis optimization
-- TODO: Test with different input sizes
--
-- ============================================================================
-- STEP 5: ADVANCED FEATURES AND OPTIMIZATIONS
-- ============================================================================
--
-- CASCADING CAPABILITY:
-- - Enable input chaining for larger encoders
-- - Priority input from higher-level encoder
-- - Group select outputs for hierarchical systems
-- - Expandable to arbitrary input counts
--
-- MASKING AND SELECTIVE ENCODING:
-- - Mask input for selective priority encoding
-- - Dynamic priority modification
-- - Conditional encoding based on system state
-- - Flexible priority assignment
--
-- MULTIPLE OUTPUT FORMATS:
-- - Binary encoded output (standard)
-- - One-hot encoded output (decoded form)
-- - Gray code encoded output (glitch reduction)
-- - BCD encoded output (decimal representation)
--
-- PERFORMANCE OPTIMIZATIONS:
-- - Parallel priority detection
-- - Carry-lookahead style encoding
-- - LUT optimization for FPGA targets
-- - Critical path minimization
--
-- TODO: Implement cascading capability
-- TODO: Add masking functionality
-- TODO: Create multiple output formats
-- TODO: Optimize for target architecture
--
-- ============================================================================
-- IMPLEMENTATION CONSIDERATIONS:
-- ============================================================================
--
-- PRIORITY ENCODING OPERATIONS:
-- - Highest priority input identification
-- - Binary position encoding
-- - Valid output generation
-- - Multiple request handling
-- - Priority conflict resolution
--
-- LOGIC OPTIMIZATION:
-- - Minimize gate count for encoding logic
-- - Optimize critical path timing
-- - Resource sharing between functions
-- - LUT utilization optimization for FPGAs
-- - Don't-care condition exploitation
--
-- TIMING CONSIDERATIONS:
-- - Propagation delay through priority logic
-- - Critical path from inputs to outputs
-- - Glitch-free operation during transitions
-- - Setup and hold time requirements
-- - Output stability during input changes
--
-- VHDL TECHNIQUES:
-- - Loop constructs for scalability
-- - Generic parameters for flexibility
-- - Type conversions for encoding
-- - Process vs. concurrent statement trade-offs
-- - Synthesis optimization attributes
--
-- SYNTHESIS CONSIDERATIONS:
-- - Priority encoder inference by tools
-- - Resource utilization (LUTs, logic elements)
-- - Critical path optimization
-- - Power consumption minimization
-- - Area vs. speed trade-offs
--
-- TESTABILITY FEATURES:
-- - Comprehensive priority pattern testing
-- - Boundary condition verification
-- - Multiple request scenario testing
-- - Random input pattern testing
-- - Built-in self-test capabilities
--
-- ============================================================================
-- APPLICATIONS:
-- ============================================================================
--
-- 1. INTERRUPT CONTROLLERS:
--    - Interrupt request prioritization
--    - Vector generation for interrupt service
--    - Nested interrupt handling
--    - Interrupt masking and control
--    - Real-time system interrupt management
--
-- 2. ARBITRATION CIRCUITS:
--    - Bus arbitration for multiple masters
--    - Resource allocation in multiprocessor systems
--    - Memory access arbitration
--    - I/O device access control
--    - Network packet scheduling
--
-- 3. PROCESSOR CONTROL UNITS:
--    - Instruction priority handling
--    - Exception and trap prioritization
--    - Pipeline hazard resolution
--    - Branch prediction priority
--    - Cache miss handling priority
--
-- 4. COMMUNICATION SYSTEMS:
--    - Message queue priority handling
--    - Protocol layer prioritization
--    - Quality of Service (QoS) implementation
--    - Traffic shaping and scheduling
--    - Error handling prioritization
--
-- 5. REAL-TIME SYSTEMS:
--    - Task scheduling priority encoding
--    - Event priority management
--    - Resource contention resolution
--    - Deadline-driven scheduling
--    - Critical section access control
--
-- 6. DIGITAL SIGNAL PROCESSING:
--    - Sample priority in multi-channel systems
--    - Filter coefficient selection
--    - Algorithm priority switching
--    - Data path selection
--    - Processing resource allocation
--
-- ============================================================================
-- TESTING STRATEGY:
-- ============================================================================
--
-- FUNCTIONAL TESTING:
-- - Test all single input activations
-- - Verify priority ordering correctness
-- - Test multiple simultaneous inputs
-- - Validate encoding accuracy
-- - Check valid output generation
--
-- PRIORITY TESTING:
-- - Highest priority input verification
-- - Lower priority input masking
-- - Priority conflict resolution
-- - Edge case priority handling
-- - Dynamic priority changes
--
-- BOUNDARY TESTING:
-- - All inputs inactive (no request)
-- - All inputs active (maximum conflict)
-- - Single input patterns
-- - Adjacent priority conflicts
-- - Wraparound conditions
--
-- ENABLE CONTROL TESTING:
-- - Enable/disable functionality
-- - Output behavior when disabled
-- - Enable timing relationships
-- - Glitch-free enable transitions
-- - Power-down mode behavior
--
-- PERFORMANCE TESTING:
-- - Propagation delay measurement
-- - Critical path identification
-- - Resource utilization analysis
-- - Power consumption measurement
-- - Temperature and voltage testing
--
-- INTEGRATION TESTING:
-- - Interrupt controller integration
-- - Arbitration system integration
-- - Processor control unit integration
-- - System-level functionality testing
-- - Multi-encoder coordination
--
-- ============================================================================
-- RECOMMENDED IMPLEMENTATION APPROACH:
-- ============================================================================
--
-- FOR BEGINNERS:
-- 1. Start with behavioral architecture using if-then-elsif
-- 2. Implement basic 4-input or 8-input encoder
-- 3. Add enable control functionality
-- 4. Create simple testbench for basic functionality
-- 5. Verify with known priority scenarios
--
-- FOR INTERMEDIATE USERS:
-- 1. Implement complete priority encoding with all features
-- 2. Add cascading capability for larger inputs
-- 3. Create comprehensive testbench with edge cases
-- 4. Analyze timing and resource utilization
-- 5. Compare different architectural approaches
--
-- FOR ADVANCED USERS:
-- 1. Implement optimized loop-based parameterized design
-- 2. Create hierarchical scalable architecture
-- 3. Optimize for specific FPGA architectures
-- 4. Implement advanced features (masking, multiple formats)
-- 5. Create reusable priority encoder library
--
-- ============================================================================
-- EXTENSION EXERCISES:
-- ============================================================================
--
-- 1. PARAMETERIZED PRIORITY ENCODER:
--    - Create generic design for any input count
--    - Implement automatic output width calculation
--    - Add compile-time priority direction selection
--    - Support runtime priority reconfiguration
--
-- 2. ROTATING PRIORITY ENCODER:
--    - Implement round-robin priority rotation
--    - Add fairness mechanisms
--    - Create aging-based priority adjustment
--    - Implement weighted priority schemes
--
-- 3. MULTI-LEVEL PRIORITY ENCODER:
--    - Implement hierarchical priority levels
--    - Add group-based priority encoding
--    - Create nested priority structures
--    - Support priority inheritance mechanisms
--
-- 4. MASKED PRIORITY ENCODER:
--    - Add dynamic input masking capability
--    - Implement selective priority encoding
--    - Create conditional priority assignment
--    - Add runtime mask configuration
--
-- 5. PIPELINE PRIORITY ENCODER:
--    - Create multi-stage pipeline for high frequency
--    - Add pipeline registers and control
--    - Implement hazard detection and handling
--    - Optimize pipeline for throughput
--
-- 6. CONTENT-ADDRESSABLE PRIORITY ENCODER:
--    - Combine with CAM functionality
--    - Add pattern matching with priority
--    - Implement associative priority lookup
--    - Create high-speed search with priority
--
-- ============================================================================
-- COMMON MISTAKES TO AVOID:
-- ============================================================================
--
-- 1. PRIORITY ORDER CONFUSION:
--    - Clearly define MSB vs. LSB priority convention
--    - Verify priority ordering in implementation
--    - Test priority resolution thoroughly
--    - Document priority convention clearly
--
-- 2. INCOMPLETE CASE COVERAGE:
--    - Handle all possible input combinations
--    - Ensure all outputs are driven in all cases
--    - Avoid inference of unwanted latches
--    - Check for undefined output states
--
-- 3. SYNTHESIS OPTIMIZATION PROBLEMS:
--    - Verify synthesis tool interpretation
--    - Check for combinational loops
--    - Ensure proper resource utilization
--    - Validate timing closure
--
-- 4. ENABLE CONTROL ERRORS:
--    - Implement proper enable gating
--    - Verify disabled state behavior
--    - Check for glitches during enable transitions
--    - Test enable timing relationships
--
-- 5. TESTBENCH INADEQUACY:
--    - Test all priority combinations
--    - Include comprehensive edge cases
--    - Verify timing relationships
--    - Check for output glitches
--
-- 6. SCALABILITY ISSUES:
--    - Design for easy expansion
--    - Use generic parameters appropriately
--    - Test with different input sizes
--    - Verify hierarchical composition
--
-- ============================================================================
-- DESIGN VERIFICATION CHECKLIST:
-- ============================================================================
--
-- □ Entity declaration includes all required ports
-- □ Priority ordering is clearly defined and documented
-- □ Encoding logic correctly identifies highest priority
-- □ Valid output accurately indicates active inputs
-- □ Enable control functions properly
-- □ All input combinations produce correct outputs
-- □ No unwanted latches are inferred
-- □ Timing requirements satisfied for target frequency
-- □ Synthesis results meet resource constraints
-- □ Code follows project VHDL style guidelines
-- □ Testbench provides comprehensive priority coverage
-- □ Documentation clearly explains priority convention
-- □ Signal assignments avoid combinational loops
-- □ All outputs are properly driven in all conditions
-- □ Design is scalable for different input counts
-- □ Performance meets or exceeds specifications
-- □ Power consumption is within acceptable limits
--
-- ============================================================================
-- DIGITAL DESIGN CONTEXT:
-- ============================================================================
--
-- PROCESSOR ARCHITECTURE INTEGRATION:
-- - Interrupt controller component
-- - Exception handling priority
-- - Instruction pipeline arbitration
-- - Cache miss priority handling
-- - Branch prediction priority
--
-- SYSTEM-ON-CHIP APPLICATIONS:
-- - Bus arbitration controllers
-- - Memory access prioritization
-- - I/O device scheduling
-- - Power management priority
-- - Clock domain crossing priority
--
-- PERFORMANCE METRICS:
-- - Encoding operations per second throughput
-- - Propagation delay (critical path)
-- - Area utilization (LUTs, logic elements)
-- - Power consumption (static, dynamic)
-- - Maximum operating frequency
--
-- DESIGN TRADE-OFFS:
-- - Speed vs. area utilization
-- - Functionality vs. complexity
-- - Power consumption vs. performance
-- - Flexibility vs. optimization
-- - Scalability vs. resource usage
--
-- ============================================================================
-- PHYSICAL IMPLEMENTATION NOTES:
-- ============================================================================
--
-- FPGA RESOURCE UTILIZATION:
-- - Logic Elements: ~5-15 LUTs for 8-input encoder
-- - Routing: Moderate for priority logic
-- - Registers: None required for combinational implementation
-- - Memory: None required for basic encoder
-- - DSP Blocks: Not typically used
--
-- TIMING CHARACTERISTICS:
-- - Combinational Delay: ~1-3ns for 8-input encoder
-- - Critical Path: Through priority detection logic
-- - Setup Time: Input signal requirements
-- - Hold Time: Input signal stability
-- - Clock-to-Output: For registered implementations
--
-- POWER CONSUMPTION:
-- - Static Power: FPGA leakage current
-- - Dynamic Power: Input switching activity dependent
-- - Encoding Power: Low for priority logic
-- - I/O Power: Interface signal switching
-- - Total Power: Function of utilization and frequency
--
-- DESIGN CONSTRAINTS:
-- - Timing constraints for critical paths
-- - Area constraints for resource utilization
-- - Power constraints for thermal management
-- - I/O constraints for interface compatibility
-- - Performance constraints for system requirements
--
-- ============================================================================
-- ADVANCED PRIORITY ENCODER CONCEPTS:
-- ============================================================================
--
-- HIERARCHICAL PRIORITY STRUCTURES:
-- - Multi-level priority encoding
-- - Group-based priority assignment
-- - Nested priority resolution
-- - Scalable priority architectures
-- - Distributed priority management
--
-- DYNAMIC PRIORITY MECHANISMS:
-- - Runtime priority reconfiguration
-- - Adaptive priority adjustment
-- - Aging-based priority modification
-- - Load-balancing priority schemes
-- - Fairness enforcement mechanisms
--
-- SPECIALIZED ENCODING TECHNIQUES:
-- - Thermometer code encoding
-- - Gray code priority encoding
-- - Weighted priority encoding
-- - Probabilistic priority selection
-- - Fuzzy priority resolution
--
-- FAULT-TOLERANT PRIORITY ENCODING:
-- - Error detection in priority logic
-- - Redundant priority encoders
-- - Graceful degradation mechanisms
-- - Self-healing priority systems
-- - Reliability enhancement techniques
--
-- ============================================================================
-- SIMULATION AND VERIFICATION NOTES:
-- ============================================================================
--
-- TESTBENCH ARCHITECTURE:
-- - Comprehensive input pattern generation
-- - Expected result calculation and comparison
-- - Priority scenario verification
-- - Edge case testing
-- - Coverage analysis and reporting
--
-- VERIFICATION METHODOLOGY:
-- - Directed testing for specific priority cases
-- - Random testing for broad coverage
-- - Constrained random testing for edge cases
-- - Formal verification for priority properties
-- - Assertion-based verification for continuous checking
--
-- DEBUGGING TECHNIQUES:
-- - Waveform analysis for priority behavior
-- - Breakpoint debugging in simulation
-- - Signal tracing through priority logic
-- - Priority conflict analysis
-- - Performance bottleneck identification
--
-- PERFORMANCE ANALYSIS:
-- - Priority encoding timing characterization
-- - Critical path identification and optimization
-- - Resource utilization vs. performance trade-offs
-- - Power analysis for different input patterns
-- - Scalability analysis for larger input counts
--
-- ============================================================================
-- IMPLEMENTATION TEMPLATE:
-- ============================================================================
--
-- [Add your library declarations here]
--
-- [Add your entity declaration here]
--
-- [Add your architecture implementation here]
--
-- ============================================================================