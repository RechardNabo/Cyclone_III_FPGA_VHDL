-- ============================================================================
-- 4-Bit Counter Implementation - Programming Guidance
-- ============================================================================
-- 
-- PROJECT OVERVIEW:
-- This file implements a 4-bit binary counter, a fundamental sequential logic
-- circuit that counts from 0 to 15 (or other ranges) in binary. Counters are
-- essential components in digital systems for timing, addressing, frequency
-- division, and control applications. They can be implemented as synchronous
-- or asynchronous designs with various counting modes and control features.
--
-- LEARNING OBJECTIVES:
-- 1. Understand sequential logic design principles
-- 2. Learn synchronous vs asynchronous counter design
-- 3. Practice clocked process implementation in VHDL
-- 4. Explore different counting modes (up, down, up/down)
-- 5. Understand counter control signals (enable, reset, load)
--
-- ============================================================================
-- STEP-BY-STEP IMPLEMENTATION GUIDE:
-- ============================================================================
--
-- STEP 1: LIBRARY DECLARATIONS
-- ----------------------------------------------------------------------------
-- Required Libraries:
-- - IEEE library for standard logic types
-- - std_logic_1164 package for std_logic and logical operators
-- - numeric_std package for arithmetic operations (recommended)
-- - std_logic_arith and std_logic_unsigned (alternative, not recommended)
-- 
-- TODO: Add library IEEE;
-- TODO: Add use IEEE.std_logic_1164.all;
-- TODO: Add use IEEE.numeric_std.all; (recommended approach)
-- TODO: Consider use IEEE.std_logic_arith.all; (alternative approach)
--
-- ============================================================================
-- STEP 2: ENTITY DECLARATION
-- ============================================================================
-- The entity defines the interface for the 4-bit counter
--
-- Entity Requirements:
-- - Name: counter_4bit (maintain current naming convention)
-- - Inputs: Clock, reset, enable, load, direction control
-- - Outputs: 4-bit count value, terminal count flags
-- - Consider different counting modes and control options
--
-- Port Specifications:
-- - clk : in std_logic (Clock input for synchronous operation)
-- - reset : in std_logic (Asynchronous or synchronous reset)
-- - enable : in std_logic (Count enable control)
-- - load : in std_logic (Parallel load control)
-- - up_down : in std_logic (Count direction: '1' = up, '0' = down)
-- - load_data : in std_logic_vector(3 downto 0) (Parallel load data)
-- - count : out std_logic_vector(3 downto 0) (Current count value)
-- - tc_up : out std_logic (Terminal count up flag - count = 15)
-- - tc_down : out std_logic (Terminal count down flag - count = 0)
-- - carry_out : out std_logic (Carry output for cascading)
-- - borrow_out : out std_logic (Borrow output for cascading)
--
-- Design Considerations:
-- - Reset type: asynchronous vs synchronous
-- - Enable type: count enable vs clock enable
-- - Load priority vs count priority
-- - Terminal count detection logic
--
-- TODO: Declare entity with appropriate port names
-- TODO: Add detailed port comments
-- TODO: Consider different control signal combinations
-- TODO: Plan for cascading capability
--
-- ============================================================================
-- STEP 3: COUNTER OPERATION DEFINITIONS
-- ============================================================================
--
-- COUNTER PRINCIPLES:
-- - Sequential logic with memory (flip-flops)
-- - State transitions on clock edges
-- - Binary counting sequence: 0, 1, 2, ..., 15, 0, ...
-- - Control signals modify counting behavior
-- - Terminal count detection for overflow/underflow
--
-- COUNTING MODES:
-- 1. UP COUNTER: 0 → 1 → 2 → ... → 15 → 0 (with wraparound)
-- 2. DOWN COUNTER: 15 → 14 → 13 → ... → 0 → 15 (with wraparound)
-- 3. UP/DOWN COUNTER: Direction controlled by up_down signal
-- 4. MODULO-N COUNTER: Count to specific value then reset
--
-- CONTROL SIGNAL BEHAVIOR:
-- - RESET: Initialize counter to 0 (or preset value)
-- - ENABLE: Allow/prevent counting operation
-- - LOAD: Parallel load of data into counter
-- - UP_DOWN: Select counting direction
--
-- PRIORITY HIERARCHY (typical):
-- 1. RESET (highest priority)
-- 2. LOAD (parallel load)
-- 3. ENABLE + UP_DOWN (counting)
-- 4. HOLD (no change when disabled)
--
-- TERMINAL COUNT CONDITIONS:
-- - TC_UP: count = "1111" (15) for up counting
-- - TC_DOWN: count = "0000" (0) for down counting
-- - Used for cascading multiple counters
-- - Can trigger external events or interrupts
--
-- TODO: Define counting state transitions
-- TODO: Plan control signal priority
-- TODO: Design terminal count logic
-- TODO: Consider edge cases and boundary conditions
--
-- ============================================================================
-- STEP 4: ARCHITECTURE IMPLEMENTATION OPTIONS
-- ============================================================================
--
-- OPTION 1: SYNCHRONOUS BEHAVIORAL ARCHITECTURE
-- ----------------------------------------------------------------------------
-- Use clocked process with synchronous design principles
--
-- Implementation Approach:
-- - Single clocked process for all sequential logic
-- - Synchronous reset and control signals
-- - Use unsigned type for arithmetic operations
-- - Clean, predictable timing behavior
--
-- Example Structure:
-- architecture behavioral of counter_4bit is
--     signal count_reg : unsigned(3 downto 0) := (others => '0');
-- begin
--     -- Main counter process
--     counter_process: process(clk)
--     begin
--         if rising_edge(clk) then
--             if reset = '1' then
--                 count_reg <= (others => '0');
--             elsif load = '1' then
--                 count_reg <= unsigned(load_data);
--             elsif enable = '1' then
--                 if up_down = '1' then
--                     count_reg <= count_reg + 1;
--                 else
--                     count_reg <= count_reg - 1;
--                 end if;
--             end if;
--         end if;
--     end process;
--     
--     -- Output assignments
--     count <= std_logic_vector(count_reg);
--     tc_up <= '1' when count_reg = 15 else '0';
--     tc_down <= '1' when count_reg = 0 else '0';
--     carry_out <= tc_up and enable and up_down;
--     borrow_out <= tc_down and enable and not up_down;
-- end behavioral;
--
-- TODO: Implement synchronous clocked process
-- TODO: Add proper reset handling
-- TODO: Implement load and enable logic
-- TODO: Generate terminal count flags
--
-- OPTION 2: ASYNCHRONOUS RESET ARCHITECTURE
-- ----------------------------------------------------------------------------
-- Use asynchronous reset for immediate counter initialization
--
-- Implementation Approach:
-- - Asynchronous reset in process sensitivity list
-- - Immediate reset response independent of clock
-- - Synchronous operation for all other controls
-- - Common in systems requiring immediate reset
--
-- Example Structure:
-- counter_process: process(clk, reset)
-- begin
--     if reset = '1' then
--         count_reg <= (others => '0');
--     elsif rising_edge(clk) then
--         if load = '1' then
--             count_reg <= unsigned(load_data);
--         elsif enable = '1' then
--             if up_down = '1' then
--                 count_reg <= count_reg + 1;
--             else
--                 count_reg <= count_reg - 1;
--             end if;
--         end if;
--     end if;
-- end process;
--
-- TODO: Implement asynchronous reset logic
-- TODO: Ensure proper reset timing
-- TODO: Verify reset priority over other controls
-- TODO: Test reset behavior in simulation
--
-- OPTION 3: MODULAR COUNTER ARCHITECTURE
-- ----------------------------------------------------------------------------
-- Implement configurable modulo-N counting
--
-- Implementation Approach:
-- - Add modulus parameter or input
-- - Reset counter when reaching modulus value
-- - Flexible counting range configuration
-- - Useful for frequency division applications
--
-- Example Structure:
-- architecture modular of counter_4bit is
--     signal count_reg : unsigned(3 downto 0) := (others => '0');
--     constant MODULUS : integer := 10; -- Count 0 to 9
-- begin
--     counter_process: process(clk, reset)
--     begin
--         if reset = '1' then
--             count_reg <= (others => '0');
--         elsif rising_edge(clk) then
--             if load = '1' then
--                 count_reg <= unsigned(load_data);
--             elsif enable = '1' then
--                 if up_down = '1' then
--                     if count_reg = MODULUS - 1 then
--                         count_reg <= (others => '0');
--                     else
--                         count_reg <= count_reg + 1;
--                     end if;
--                 else
--                     if count_reg = 0 then
--                         count_reg <= to_unsigned(MODULUS - 1, 4);
--                     else
--                         count_reg <= count_reg - 1;
--                     end if;
--                 end if;
--             end if;
--         end if;
--     end process;
-- end modular;
--
-- TODO: Implement modulus parameter
-- TODO: Add modulo counting logic
-- TODO: Update terminal count conditions
-- TODO: Test different modulus values
--
-- OPTION 4: CASCADABLE COUNTER ARCHITECTURE
-- ----------------------------------------------------------------------------
-- Design for easy cascading with other counters
--
-- Implementation Approach:
-- - Add carry/borrow inputs and outputs
-- - Enable cascading for wider counters
-- - Proper terminal count generation
-- - Chain multiple 4-bit counters
--
-- Example Structure:
-- entity counter_4bit is
--     port (
--         clk : in std_logic;
--         reset : in std_logic;
--         enable : in std_logic;
--         carry_in : in std_logic;
--         borrow_in : in std_logic;
--         up_down : in std_logic;
--         count : out std_logic_vector(3 downto 0);
--         carry_out : out std_logic;
--         borrow_out : out std_logic
--     );
-- end counter_4bit;
--
-- -- Enable logic for cascading
-- enable_internal <= enable and ((carry_in and up_down) or (borrow_in and not up_down));
--
-- TODO: Add cascade input/output ports
-- TODO: Implement cascade enable logic
-- TODO: Generate proper carry/borrow signals
-- TODO: Test cascaded counter operation
--
-- ============================================================================
-- STEP 5: ADVANCED COUNTER FEATURES
-- ============================================================================
--
-- PRESET COUNTER:
-- - Initialize to specific value instead of zero
-- - Useful for countdown timers
-- - Configurable preset value
-- - Preset enable control signal
--
-- GRAY CODE COUNTER:
-- - Only one bit changes per count
-- - Reduces switching noise and power
-- - Useful for asynchronous interfaces
-- - Requires Gray code conversion logic
--
-- JOHNSON COUNTER (RING COUNTER):
-- - Shift register with inverted feedback
-- - 2N states for N flip-flops
-- - Self-starting with proper initialization
-- - Useful for timing and control sequences
--
-- BCD COUNTER:
-- - Binary Coded Decimal counting (0-9)
-- - Reset at count 10 instead of 16
-- - Useful for decimal displays
-- - Multiple BCD digits for larger numbers
--
-- PROGRAMMABLE COUNTER:
-- - Runtime configurable count sequence
-- - Load different modulus values
-- - Flexible timing generation
-- - Microprocessor-controlled operation
--
-- TODO: Choose appropriate advanced features
-- TODO: Implement selected counter type
-- TODO: Add necessary control logic
-- TODO: Verify advanced functionality
--
-- ============================================================================
-- IMPLEMENTATION CONSIDERATIONS:
-- ============================================================================
--
-- SEQUENTIAL LOGIC DESIGN:
-- - Proper clocking methodology
-- - Setup and hold time requirements
-- - Clock domain considerations
-- - Reset strategy (sync vs async)
-- - Metastability prevention
--
-- TIMING CONSIDERATIONS:
-- - Clock-to-output delay
-- - Setup time for control signals
-- - Hold time requirements
-- - Clock skew tolerance
-- - Maximum operating frequency
--
-- VHDL TECHNIQUES:
-- - Process sensitivity lists
-- - Signal vs variable usage
-- - Type conversions (std_logic_vector ↔ unsigned)
-- - Concurrent vs sequential statements
-- - Synthesis optimization attributes
--
-- SYNTHESIS CONSIDERATIONS:
-- - Flip-flop inference
-- - Resource utilization optimization
-- - Clock domain crossing
-- - Reset tree optimization
-- - Power optimization techniques
--
-- TESTABILITY FEATURES:
-- - Comprehensive test patterns
-- - Boundary condition testing
-- - Control signal interaction testing
-- - Timing verification
-- - Built-in self-test capabilities
--
-- ============================================================================
-- APPLICATIONS:
-- ============================================================================
--
-- 1. FREQUENCY DIVISION:
--    - Clock frequency reduction
--    - Timing signal generation
--    - Baud rate generation for UARTs
--    - PWM frequency control
--    - System clock derivation
--
-- 2. ADDRESS GENERATION:
--    - Memory address counters
--    - ROM/RAM addressing
--    - Sequential memory access
--    - DMA address generation
--    - Cache line addressing
--
-- 3. TIMING AND CONTROL:
--    - State machine timing
--    - Delay generation
--    - Timeout counters
--    - Watchdog timers
--    - Event counting
--
-- 4. DIGITAL DISPLAYS:
--    - 7-segment display control
--    - LED matrix scanning
--    - Multiplexed display timing
--    - Digit selection control
--    - Display refresh timing
--
-- 5. COMMUNICATION PROTOCOLS:
--    - Bit counting in serial protocols
--    - Frame counting
--    - Packet sequence numbers
--    - Protocol timeout handling
--    - Error retry counting
--
-- 6. SIGNAL PROCESSING:
--    - Sample counting
--    - Window function control
--    - Filter coefficient indexing
--    - FFT butterfly control
--    - Decimation and interpolation
--
-- ============================================================================
-- TESTING STRATEGY:
-- ============================================================================
--
-- FUNCTIONAL TESTING:
-- - Test complete count sequence (0 to 15)
-- - Verify wraparound behavior
-- - Test up and down counting modes
-- - Validate control signal functionality
-- - Check terminal count flag generation
--
-- CONTROL SIGNAL TESTING:
-- - Reset functionality (sync/async)
-- - Enable control behavior
-- - Load operation verification
-- - Up/down direction control
-- - Control signal priority testing
--
-- BOUNDARY CONDITION TESTING:
-- - Count overflow (15 → 0)
-- - Count underflow (0 → 15)
-- - Maximum count value behavior
-- - Minimum count value behavior
-- - Edge case combinations
--
-- TIMING TESTING:
-- - Setup and hold time verification
-- - Clock edge sensitivity
-- - Propagation delay measurement
-- - Control signal timing relationships
-- - Metastability testing
--
-- INTEGRATION TESTING:
-- - Cascaded counter operation
-- - System-level integration
-- - Clock domain crossing
-- - Reset distribution testing
-- - Performance under load
--
-- ============================================================================
-- RECOMMENDED IMPLEMENTATION APPROACH:
-- ============================================================================
--
-- FOR BEGINNERS:
-- 1. Start with simple synchronous up counter
-- 2. Add basic reset functionality
-- 3. Implement enable control
-- 4. Create simple testbench
-- 5. Verify basic counting operation
--
-- FOR INTERMEDIATE USERS:
-- 1. Add up/down counting capability
-- 2. Implement parallel load feature
-- 3. Add terminal count flag generation
-- 4. Create comprehensive testbench
-- 5. Analyze timing and resource usage
--
-- FOR ADVANCED USERS:
-- 1. Implement cascadable counter design
-- 2. Add advanced features (preset, modulo)
-- 3. Optimize for specific FPGA architecture
-- 4. Create parameterized generic design
-- 5. Implement built-in self-test features
--
-- ============================================================================
-- EXTENSION EXERCISES:
-- ============================================================================
--
-- 1. N-BIT PARAMETERIZED COUNTER:
--    - Generic bit width parameter
--    - Scalable to any size
--    - Automatic terminal count calculation
--    - Resource optimization for different sizes
--
-- 2. MULTI-MODE COUNTER:
--    - Binary, BCD, Gray code modes
--    - Runtime mode selection
--    - Mode-specific terminal counts
--    - Unified control interface
--
-- 3. PRESCALER COUNTER:
--    - Configurable prescale ratios
--    - Fractional frequency division
--    - Duty cycle control
--    - Phase alignment features
--
-- 4. COUNTER WITH INTERRUPTS:
--    - Interrupt generation on terminal count
--    - Programmable interrupt thresholds
--    - Interrupt masking and control
--    - Priority interrupt handling
--
-- 5. FAULT-TOLERANT COUNTER:
--    - Error detection and correction
--    - Redundant counting logic
--    - Self-checking capabilities
--    - Graceful degradation modes
--
-- 6. HIGH-SPEED COUNTER:
--    - Pipeline architecture for high frequency
--    - Parallel counting techniques
--    - Clock domain optimization
--    - Timing closure optimization
--
-- ============================================================================
-- COMMON MISTAKES TO AVOID:
-- ============================================================================
--
-- 1. CLOCKING ISSUES:
--    - Multiple clock edges in process
--    - Incomplete sensitivity lists
--    - Clock domain crossing problems
--    - Gated clock usage
--
-- 2. RESET PROBLEMS:
--    - Incomplete reset conditions
--    - Reset signal timing issues
--    - Mixed sync/async reset usage
--    - Reset priority conflicts
--
-- 3. CONTROL SIGNAL CONFLICTS:
--    - Undefined priority between controls
--    - Simultaneous conflicting controls
--    - Control signal setup violations
--    - Enable logic errors
--
-- 4. TYPE CONVERSION ERRORS:
--    - Incorrect std_logic_vector ↔ unsigned conversion
--    - Size mismatch in assignments
--    - Signed vs unsigned arithmetic
--    - Range check failures
--
-- 5. SYNTHESIS ISSUES:
--    - Unwanted latch inference
--    - Incomplete case statements
--    - Non-synthesizable constructs
--    - Resource utilization problems
--
-- 6. TESTBENCH INADEQUACY:
--    - Insufficient test coverage
--    - Missing edge cases
--    - Incorrect timing relationships
--    - Inadequate verification methodology
--
-- ============================================================================
-- DESIGN VERIFICATION CHECKLIST:
-- ============================================================================
--
-- □ Entity declaration includes all required ports
-- □ Clock and reset signals properly handled
-- □ Count sequence operates correctly
-- □ Control signals function as specified
-- □ Terminal count flags generated accurately
-- □ No unwanted latches inferred
-- □ Timing requirements satisfied
-- □ Synthesis results meet resource constraints
-- □ Code follows VHDL style guidelines
-- □ Testbench provides comprehensive coverage
-- □ Documentation clearly explains operation
-- □ All outputs properly driven
-- □ Design scalable for different applications
-- □ Performance meets specifications
-- □ Power consumption acceptable
--
-- ============================================================================
-- DIGITAL DESIGN CONTEXT:
-- ============================================================================
--
-- SEQUENTIAL LOGIC FUNDAMENTALS:
-- - State storage using flip-flops
-- - Clock-driven state transitions
-- - Memory elements in digital systems
-- - Synchronous design methodology
-- - Timing analysis and constraints
--
-- SYSTEM INTEGRATION:
-- - Counter as building block
-- - Interface with combinational logic
-- - Clock domain considerations
-- - Reset distribution networks
-- - Power management integration
--
-- PERFORMANCE METRICS:
-- - Maximum counting frequency
-- - Power consumption per count
-- - Resource utilization efficiency
-- - Setup/hold time margins
-- - Jitter and timing accuracy
--
-- DESIGN TRADE-OFFS:
-- - Speed vs power consumption
-- - Functionality vs complexity
-- - Area vs performance
-- - Flexibility vs optimization
-- - Testability vs efficiency
--
-- ============================================================================
-- PHYSICAL IMPLEMENTATION NOTES:
-- ============================================================================
--
-- FPGA RESOURCE UTILIZATION:
-- - Logic Elements: ~4-6 LUTs for 4-bit counter
-- - Registers: 4 flip-flops for count storage
-- - Routing: Moderate for control signals
-- - Memory: None required for basic counter
-- - Clock Resources: Global clock networks
--
-- TIMING CHARACTERISTICS:
-- - Clock-to-Output: ~1-3ns typical
-- - Setup Time: Control signal requirements
-- - Hold Time: Input signal stability
-- - Maximum Frequency: 200-500MHz typical
-- - Jitter: Clock quality dependent
--
-- POWER CONSUMPTION:
-- - Static Power: Flip-flop leakage
-- - Dynamic Power: Switching activity dependent
-- - Clock Power: Clock tree distribution
-- - I/O Power: Output signal switching
-- - Total Power: Function of frequency and activity
--
-- DESIGN CONSTRAINTS:
-- - Timing constraints for clock domains
-- - Reset timing and distribution
-- - Control signal setup/hold requirements
-- - Power consumption limits
-- - Resource utilization targets
--
-- ============================================================================
-- IMPLEMENTATION TEMPLATE:
-- ============================================================================
--
-- [Add your library declarations here]
--
-- [Add your entity declaration here]
--
-- [Add your architecture implementation here]
--
-- ============================================================================