-- Cortex-A72 Interface VHDL File
-- This file contains the interface definition for ARM Cortex-A72 processor
-- 
-- Author: [To be filled]
-- Date: [To be filled]
-- Description: Interface module for Cortex-A72 processor integration

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-- Entity declaration will be added here
-- Interface signals and ports will be defined here
-- Implementation to be completed